library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity game_rom is
    Port ( address : in STD_LOGIC_VECTOR (15 downto 0);
           clock : in STD_LOGIC;
           we : in STD_LOGIC;
           dataIn : in STD_LOGIC_VECTOR (7 downto 0);
           dataOut : out STD_LOGIC_VECTOR (7 downto 0));
end game_rom;

architecture Behavioral of game_rom is
    type RAM is array ( ( 16 * 4096 ) - 1 downto 0 ) of std_logic_vector( 7 downto 0 );
    
    signal sys_RAM : RAM := (   
                                -- light travels left
                                (0 + 136) => x"00", (0 + 137) => x"00", -- delay
                                (0 + 138) => x"00",
                                512 => x"66", 513 => x"01",  -- LD V6, 0x01
                                514 => x"61", 515 => x"3C",  -- LD V1, 0x3C
                                516 => x"F1", 517 => x"15",  -- LD DT, V1;   ; loop
                                518 => x"86", 519 => x"6E",  -- SHL V6, V6
                                520 => x"4F", 521 => x"01",  -- SNE VF, 0x01
                                522 => x"66", 523 => x"01",  -- LD V6, 0x01
                                524 => x"80", 525 => x"60",  -- LD V0, V6
                                526 => x"A1", 527 => x"FF",  -- LD I, 0x1FF
                                528 => x"F0", 529 => x"55",  -- LD [I], V0
                                530 => x"F2", 531 => x"07",  -- LD V2, DT   ; wait
                                532 => x"32", 533 => x"00",  -- SE V2, 0x00
                                534 => x"12", 535 => x"12",  -- JP wait
                                536 => x"12", 537 => x"04",  -- JP loop
                                
                                -- light travels right
                                (4096 + 136) => x"00", (4096 + 137) => x"00", -- delay
                                (4096 + 138) => x"00",
                                (4096 + 512) => x"66", (4096 + 513) => x"80",  -- LD V6, 0x80
                                (4096 + 514) => x"61", (4096 + 515) => x"3C",  -- LD V1, 0x3C
                                (4096 + 516) => x"F1", (4096 + 517) => x"15",  -- LD DT, V1;   ; loop
                                (4096 + 518) => x"86", (4096 + 519) => x"66",  -- SHR V6, V6
                                (4096 + 520) => x"4F", (4096 + 521) => x"01",  -- SNE VF, 0x01
                                (4096 + 522) => x"66", (4096 + 523) => x"80",  -- LD V6, 0x80
                                (4096 + 524) => x"80", (4096 + 525) => x"60",  -- LD V0, V6
                                (4096 + 526) => x"A1", (4096 + 527) => x"FF",  -- LD I, 0x1FF
                                (4096 + 528) => x"F0", (4096 + 529) => x"55",  -- LD [I], V0
                                (4096 + 530) => x"F2", (4096 + 531) => x"07",  -- LD V2, DT   ; wait
                                (4096 + 532) => x"32", (4096 + 533) => x"00",  -- SE V2, 0x00
                                (4096 + 534) => x"12", (4096 + 535) => x"12",  -- JP wait
                                (4096 + 536) => x"12", (4096 + 537) => x"04",  -- JP loop
                                
                                -- random lights
                                (8192 + 136) => x"00", (8192 + 137) => x"00", -- delay
                                (8192 + 138) => x"00",
                                (8192 + 512) => x"61", (8192 + 513) => x"3C",  -- LD V1, 0x3C
                                (8192 + 514) => x"F1", (8192 + 515) => x"15",  -- LD DT, V1;   ; loop
                                (8192 + 516) => x"C0", (8192 + 517) => x"FF",  -- RND V0, FF
                                (8192 + 518) => x"A1", (8192 + 519) => x"FF",  -- LD I, 0x1FF
                                (8192 + 520) => x"F0", (8192 + 521) => x"55",  -- LD [I], V0
                                (8192 + 522) => x"F2", (8192 + 523) => x"07",  -- LD V2, DT   ; wait
                                (8192 + 524) => x"32", (8192 + 525) => x"00",  -- SE V2, 0x00
                                (8192 + 526) => x"12", (8192 + 527) => x"0A",  -- JP wait
                                (8192 + 528) => x"12", (8192 + 529) => x"02",  -- JP loop
                                

                                -- PONG by Paul Vervalin
                                (12288 + 128) => x"0C", (12288 + 129) => x"00", 
                                (12288 + 130) => x"F0", (12288 + 131) => x"00",
                                (12288 + 132) => x"00", (12288 + 133) => x"00",
                                (12288 + 134) => x"BE", (12288 + 135) => x"00",
                                (12288 + 136) => x"00", (12288 + 137) => x"30", -- delay
                                (12288 + 138) => x"00",
                                (12288 + 512) => x"6a", (12288 + 513) => x"02", (12288 + 514) => x"6b", (12288 + 515) => x"0c", (12288 + 516) => x"6c", (12288 + 517) => x"3f", (12288 + 518) => x"6d", (12288 + 519) => x"0c", (12288 + 520) => x"a2", (12288 + 521) => x"ea", (12288 + 522) => x"da", (12288 + 523) => x"b6", (12288 + 524) => x"dc", (12288 + 525) => x"d6", (12288 + 526) => x"6e", (12288 + 527) => x"00", (12288 + 528) => x"22", (12288 + 529) => x"d4", (12288 + 530) => x"66", (12288 + 531) => x"03", (12288 + 532) => x"68", (12288 + 533) => x"02", (12288 + 534) => x"60", (12288 + 535) => x"60", (12288 + 536) => x"f0", (12288 + 537) => x"15", (12288 + 538) => x"f0", (12288 + 539) => x"07", (12288 + 540) => x"30", (12288 + 541) => x"00", (12288 + 542) => x"12", (12288 + 543) => x"1a", (12288 + 544) => x"c7", (12288 + 545) => x"17", (12288 + 546) => x"77", (12288 + 547) => x"08", (12288 + 548) => x"69", (12288 + 549) => x"ff", (12288 + 550) => x"a2", (12288 + 551) => x"f0", (12288 + 552) => x"d6", (12288 + 553) => x"71", (12288 + 554) => x"a2", (12288 + 555) => x"ea", (12288 + 556) => x"da", (12288 + 557) => x"b6", (12288 + 558) => x"dc", (12288 + 559) => x"d6", (12288 + 560) => x"60", (12288 + 561) => x"01", (12288 + 562) => x"e0", (12288 + 563) => x"a1", (12288 + 564) => x"7b", (12288 + 565) => x"fe", (12288 + 566) => x"60", (12288 + 567) => x"04", (12288 + 568) => x"e0", (12288 + 569) => x"a1", (12288 + 570) => x"7b", (12288 + 571) => x"02", (12288 + 572) => x"60", (12288 + 573) => x"1f", (12288 + 574) => x"8b", (12288 + 575) => x"02", (12288 + 576) => x"da", (12288 + 577) => x"b6", (12288 + 578) => x"60", (12288 + 579) => x"0c", (12288 + 580) => x"e0", (12288 + 581) => x"a1", (12288 + 582) => x"7d", (12288 + 583) => x"fe", (12288 + 584) => x"60", (12288 + 585) => x"0d", (12288 + 586) => x"e0", (12288 + 587) => x"a1", (12288 + 588) => x"7d", (12288 + 589) => x"02", (12288 + 590) => x"60", (12288 + 591) => x"1f", (12288 + 592) => x"8d", (12288 + 593) => x"02", (12288 + 594) => x"dc", (12288 + 595) => x"d6", (12288 + 596) => x"a2", (12288 + 597) => x"f0", (12288 + 598) => x"d6", (12288 + 599) => x"71", (12288 + 600) => x"86", (12288 + 601) => x"84", (12288 + 602) => x"87", (12288 + 603) => x"94", (12288 + 604) => x"60", (12288 + 605) => x"3f", (12288 + 606) => x"86", (12288 + 607) => x"02", (12288 + 608) => x"61", (12288 + 609) => x"1f", (12288 + 610) => x"87", (12288 + 611) => x"12", (12288 + 612) => x"46", (12288 + 613) => x"02", (12288 + 614) => x"12", (12288 + 615) => x"78", (12288 + 616) => x"46", (12288 + 617) => x"3f", (12288 + 618) => x"12", (12288 + 619) => x"82", (12288 + 620) => x"47", (12288 + 621) => x"1f", (12288 + 622) => x"69", (12288 + 623) => x"ff", (12288 + 624) => x"47", (12288 + 625) => x"00", (12288 + 626) => x"69", (12288 + 627) => x"01", (12288 + 628) => x"d6", (12288 + 629) => x"71", (12288 + 630) => x"12", (12288 + 631) => x"2a", (12288 + 632) => x"68", (12288 + 633) => x"02", (12288 + 634) => x"63", (12288 + 635) => x"01", (12288 + 636) => x"80", (12288 + 637) => x"70", (12288 + 638) => x"80", (12288 + 639) => x"b5", (12288 + 640) => x"12", (12288 + 641) => x"8a", (12288 + 642) => x"68", (12288 + 643) => x"fe", (12288 + 644) => x"63", (12288 + 645) => x"0a", (12288 + 646) => x"80", (12288 + 647) => x"70", (12288 + 648) => x"80", (12288 + 649) => x"d5", (12288 + 650) => x"3f", (12288 + 651) => x"01", (12288 + 652) => x"12", (12288 + 653) => x"a2", (12288 + 654) => x"61", (12288 + 655) => x"02", (12288 + 656) => x"80", (12288 + 657) => x"15", (12288 + 658) => x"3f", (12288 + 659) => x"01", (12288 + 660) => x"12", (12288 + 661) => x"ba", (12288 + 662) => x"80", (12288 + 663) => x"15", (12288 + 664) => x"3f", (12288 + 665) => x"01", (12288 + 666) => x"12", (12288 + 667) => x"c8", (12288 + 668) => x"80", (12288 + 669) => x"15", (12288 + 670) => x"3f", (12288 + 671) => x"01", (12288 + 672) => x"12", (12288 + 673) => x"c2", (12288 + 674) => x"60", (12288 + 675) => x"20", (12288 + 676) => x"f0", (12288 + 677) => x"18", (12288 + 678) => x"22", (12288 + 679) => x"d4", (12288 + 680) => x"8e", (12288 + 681) => x"34", (12288 + 682) => x"22", (12288 + 683) => x"d4", (12288 + 684) => x"66", (12288 + 685) => x"3e", (12288 + 686) => x"33", (12288 + 687) => x"01", (12288 + 688) => x"66", (12288 + 689) => x"03", (12288 + 690) => x"68", (12288 + 691) => x"fe", (12288 + 692) => x"33", (12288 + 693) => x"01", (12288 + 694) => x"68", (12288 + 695) => x"02", (12288 + 696) => x"12", (12288 + 697) => x"16", (12288 + 698) => x"79", (12288 + 699) => x"ff", (12288 + 700) => x"49", (12288 + 701) => x"fe", (12288 + 702) => x"69", (12288 + 703) => x"ff", (12288 + 704) => x"12", (12288 + 705) => x"c8", (12288 + 706) => x"79", (12288 + 707) => x"01", (12288 + 708) => x"49", (12288 + 709) => x"02", (12288 + 710) => x"69", (12288 + 711) => x"01", (12288 + 712) => x"60", (12288 + 713) => x"04", (12288 + 714) => x"f0", (12288 + 715) => x"18", (12288 + 716) => x"76", (12288 + 717) => x"01", (12288 + 718) => x"46", (12288 + 719) => x"40", (12288 + 720) => x"76", (12288 + 721) => x"fe", (12288 + 722) => x"12", (12288 + 723) => x"6c", (12288 + 724) => x"a2", (12288 + 725) => x"f2", (12288 + 726) => x"fe", (12288 + 727) => x"33", (12288 + 728) => x"f2", (12288 + 729) => x"65", (12288 + 730) => x"f1", (12288 + 731) => x"29", (12288 + 732) => x"64", (12288 + 733) => x"14", (12288 + 734) => x"65", (12288 + 735) => x"00", (12288 + 736) => x"d4", (12288 + 737) => x"55", (12288 + 738) => x"74", (12288 + 739) => x"15", (12288 + 740) => x"f2", (12288 + 741) => x"29", (12288 + 742) => x"d4", (12288 + 743) => x"55", (12288 + 744) => x"00", (12288 + 745) => x"ee", (12288 + 746) => x"80", (12288 + 747) => x"80", (12288 + 748) => x"80", (12288 + 749) => x"80", (12288 + 750) => x"80", (12288 + 751) => x"80", (12288 + 752) => x"80", (12288 + 753) => x"00", (12288 + 754) => x"00", (12288 + 755) => x"00", (12288 + 756) => x"00", (12288 + 757) => x"00", 
                                
                                -- Tetris by Fran Dachille
                                (16384 + 128) => x"00", (16384 + 129) => x"F0", 
                                (16384 + 130) => x"DC", (16384 + 131) => x"E0",
                                (16384 + 132) => x"F0", (16384 + 133) => x"00",
                                (16384 + 134) => x"BE", (16384 + 135) => x"00",
                                (16384 + 136) => x"00", (16384 + 137) => x"20", -- delay
                                (16384 + 138) => x"00",
                                (16384 + 512) => x"a2", (16384 + 513) => x"b4", (16384 + 514) => x"23", (16384 + 515) => x"e6", (16384 + 516) => x"22", (16384 + 517) => x"b6", (16384 + 518) => x"70", (16384 + 519) => x"01", (16384 + 520) => x"d0", (16384 + 521) => x"11", (16384 + 522) => x"30", (16384 + 523) => x"25", (16384 + 524) => x"12", (16384 + 525) => x"06", (16384 + 526) => x"71", (16384 + 527) => x"ff", (16384 + 528) => x"d0", (16384 + 529) => x"11", (16384 + 530) => x"60", (16384 + 531) => x"1a", (16384 + 532) => x"d0", (16384 + 533) => x"11", (16384 + 534) => x"60", (16384 + 535) => x"25", (16384 + 536) => x"31", (16384 + 537) => x"00", (16384 + 538) => x"12", (16384 + 539) => x"0e", (16384 + 540) => x"c4", (16384 + 541) => x"70", (16384 + 542) => x"44", (16384 + 543) => x"70", (16384 + 544) => x"12", (16384 + 545) => x"1c", (16384 + 546) => x"c3", (16384 + 547) => x"03", (16384 + 548) => x"60", (16384 + 549) => x"1e", (16384 + 550) => x"61", (16384 + 551) => x"03", (16384 + 552) => x"22", (16384 + 553) => x"5c", (16384 + 554) => x"f5", (16384 + 555) => x"15", (16384 + 556) => x"d0", (16384 + 557) => x"14", (16384 + 558) => x"3f", (16384 + 559) => x"01", (16384 + 560) => x"12", (16384 + 561) => x"3c", (16384 + 562) => x"d0", (16384 + 563) => x"14", (16384 + 564) => x"71", (16384 + 565) => x"ff", (16384 + 566) => x"d0", (16384 + 567) => x"14", (16384 + 568) => x"23", (16384 + 569) => x"40", (16384 + 570) => x"12", (16384 + 571) => x"1c", (16384 + 572) => x"e7", (16384 + 573) => x"a1", (16384 + 574) => x"22", (16384 + 575) => x"72", (16384 + 576) => x"e8", (16384 + 577) => x"a1", (16384 + 578) => x"22", (16384 + 579) => x"84", (16384 + 580) => x"e9", (16384 + 581) => x"a1", (16384 + 582) => x"22", (16384 + 583) => x"96", (16384 + 584) => x"e2", (16384 + 585) => x"9e", (16384 + 586) => x"12", (16384 + 587) => x"50", (16384 + 588) => x"66", (16384 + 589) => x"00", (16384 + 590) => x"f6", (16384 + 591) => x"15", (16384 + 592) => x"f6", (16384 + 593) => x"07", (16384 + 594) => x"36", (16384 + 595) => x"00", (16384 + 596) => x"12", (16384 + 597) => x"3c", (16384 + 598) => x"d0", (16384 + 599) => x"14", (16384 + 600) => x"71", (16384 + 601) => x"01", (16384 + 602) => x"12", (16384 + 603) => x"2a", (16384 + 604) => x"a2", (16384 + 605) => x"c4", (16384 + 606) => x"f4", (16384 + 607) => x"1e", (16384 + 608) => x"66", (16384 + 609) => x"00", (16384 + 610) => x"43", (16384 + 611) => x"01", (16384 + 612) => x"66", (16384 + 613) => x"04", (16384 + 614) => x"43", (16384 + 615) => x"02", (16384 + 616) => x"66", (16384 + 617) => x"08", (16384 + 618) => x"43", (16384 + 619) => x"03", (16384 + 620) => x"66", (16384 + 621) => x"0c", (16384 + 622) => x"f6", (16384 + 623) => x"1e", (16384 + 624) => x"00", (16384 + 625) => x"ee", (16384 + 626) => x"d0", (16384 + 627) => x"14", (16384 + 628) => x"70", (16384 + 629) => x"ff", (16384 + 630) => x"23", (16384 + 631) => x"34", (16384 + 632) => x"3f", (16384 + 633) => x"01", (16384 + 634) => x"00", (16384 + 635) => x"ee", (16384 + 636) => x"d0", (16384 + 637) => x"14", (16384 + 638) => x"70", (16384 + 639) => x"01", (16384 + 640) => x"23", (16384 + 641) => x"34", (16384 + 642) => x"00", (16384 + 643) => x"ee", (16384 + 644) => x"d0", (16384 + 645) => x"14", (16384 + 646) => x"70", (16384 + 647) => x"01", (16384 + 648) => x"23", (16384 + 649) => x"34", (16384 + 650) => x"3f", (16384 + 651) => x"01", (16384 + 652) => x"00", (16384 + 653) => x"ee", (16384 + 654) => x"d0", (16384 + 655) => x"14", (16384 + 656) => x"70", (16384 + 657) => x"ff", (16384 + 658) => x"23", (16384 + 659) => x"34", (16384 + 660) => x"00", (16384 + 661) => x"ee", (16384 + 662) => x"d0", (16384 + 663) => x"14", (16384 + 664) => x"73", (16384 + 665) => x"01", (16384 + 666) => x"43", (16384 + 667) => x"04", (16384 + 668) => x"63", (16384 + 669) => x"00", (16384 + 670) => x"22", (16384 + 671) => x"5c", (16384 + 672) => x"23", (16384 + 673) => x"34", (16384 + 674) => x"3f", (16384 + 675) => x"01", (16384 + 676) => x"00", (16384 + 677) => x"ee", (16384 + 678) => x"d0", (16384 + 679) => x"14", (16384 + 680) => x"73", (16384 + 681) => x"ff", (16384 + 682) => x"43", (16384 + 683) => x"ff", (16384 + 684) => x"63", (16384 + 685) => x"03", (16384 + 686) => x"22", (16384 + 687) => x"5c", (16384 + 688) => x"23", (16384 + 689) => x"34", (16384 + 690) => x"00", (16384 + 691) => x"ee", (16384 + 692) => x"80", (16384 + 693) => x"00", (16384 + 694) => x"67", (16384 + 695) => x"05", (16384 + 696) => x"68", (16384 + 697) => x"06", (16384 + 698) => x"69", (16384 + 699) => x"04", (16384 + 700) => x"61", (16384 + 701) => x"1f", (16384 + 702) => x"65", (16384 + 703) => x"10", (16384 + 704) => x"62", (16384 + 705) => x"07", (16384 + 706) => x"00", (16384 + 707) => x"ee", (16384 + 708) => x"40", (16384 + 709) => x"e0", (16384 + 710) => x"00", (16384 + 711) => x"00", (16384 + 712) => x"40", (16384 + 713) => x"c0", (16384 + 714) => x"40", (16384 + 715) => x"00", (16384 + 716) => x"00", (16384 + 717) => x"e0", (16384 + 718) => x"40", (16384 + 719) => x"00", (16384 + 720) => x"40", (16384 + 721) => x"60", (16384 + 722) => x"40", (16384 + 723) => x"00", (16384 + 724) => x"40", (16384 + 725) => x"40", (16384 + 726) => x"60", (16384 + 727) => x"00", (16384 + 728) => x"20", (16384 + 729) => x"e0", (16384 + 730) => x"00", (16384 + 731) => x"00", (16384 + 732) => x"c0", (16384 + 733) => x"40", (16384 + 734) => x"40", (16384 + 735) => x"00", (16384 + 736) => x"00", (16384 + 737) => x"e0", (16384 + 738) => x"80", (16384 + 739) => x"00", (16384 + 740) => x"40", (16384 + 741) => x"40", (16384 + 742) => x"c0", (16384 + 743) => x"00", (16384 + 744) => x"00", (16384 + 745) => x"e0", (16384 + 746) => x"20", (16384 + 747) => x"00", (16384 + 748) => x"60", (16384 + 749) => x"40", (16384 + 750) => x"40", (16384 + 751) => x"00", (16384 + 752) => x"80", (16384 + 753) => x"e0", (16384 + 754) => x"00", (16384 + 755) => x"00", (16384 + 756) => x"40", (16384 + 757) => x"c0", (16384 + 758) => x"80", (16384 + 759) => x"00", (16384 + 760) => x"c0", (16384 + 761) => x"60", (16384 + 762) => x"00", (16384 + 763) => x"00", (16384 + 764) => x"40", (16384 + 765) => x"c0", (16384 + 766) => x"80", (16384 + 767) => x"00", (16384 + 768) => x"c0", (16384 + 769) => x"60", (16384 + 770) => x"00", (16384 + 771) => x"00", (16384 + 772) => x"80", (16384 + 773) => x"c0", (16384 + 774) => x"40", (16384 + 775) => x"00", (16384 + 776) => x"00", (16384 + 777) => x"60", (16384 + 778) => x"c0", (16384 + 779) => x"00", (16384 + 780) => x"80", (16384 + 781) => x"c0", (16384 + 782) => x"40", (16384 + 783) => x"00", (16384 + 784) => x"00", (16384 + 785) => x"60", (16384 + 786) => x"c0", (16384 + 787) => x"00", (16384 + 788) => x"c0", (16384 + 789) => x"c0", (16384 + 790) => x"00", (16384 + 791) => x"00", (16384 + 792) => x"c0", (16384 + 793) => x"c0", (16384 + 794) => x"00", (16384 + 795) => x"00", (16384 + 796) => x"c0", (16384 + 797) => x"c0", (16384 + 798) => x"00", (16384 + 799) => x"00", (16384 + 800) => x"c0", (16384 + 801) => x"c0", (16384 + 802) => x"00", (16384 + 803) => x"00", (16384 + 804) => x"40", (16384 + 805) => x"40", (16384 + 806) => x"40", (16384 + 807) => x"40", (16384 + 808) => x"00", (16384 + 809) => x"f0", (16384 + 810) => x"00", (16384 + 811) => x"00", (16384 + 812) => x"40", (16384 + 813) => x"40", (16384 + 814) => x"40", (16384 + 815) => x"40", (16384 + 816) => x"00", (16384 + 817) => x"f0", (16384 + 818) => x"00", (16384 + 819) => x"00", (16384 + 820) => x"d0", (16384 + 821) => x"14", (16384 + 822) => x"66", (16384 + 823) => x"35", (16384 + 824) => x"76", (16384 + 825) => x"ff", (16384 + 826) => x"36", (16384 + 827) => x"00", (16384 + 828) => x"13", (16384 + 829) => x"38", (16384 + 830) => x"00", (16384 + 831) => x"ee", (16384 + 832) => x"a2", (16384 + 833) => x"b4", (16384 + 834) => x"8c", (16384 + 835) => x"10", (16384 + 836) => x"3c", (16384 + 837) => x"1e", (16384 + 838) => x"7c", (16384 + 839) => x"01", (16384 + 840) => x"3c", (16384 + 841) => x"1e", (16384 + 842) => x"7c", (16384 + 843) => x"01", (16384 + 844) => x"3c", (16384 + 845) => x"1e", (16384 + 846) => x"7c", (16384 + 847) => x"01", (16384 + 848) => x"23", (16384 + 849) => x"5e", (16384 + 850) => x"4b", (16384 + 851) => x"0a", (16384 + 852) => x"23", (16384 + 853) => x"72", (16384 + 854) => x"91", (16384 + 855) => x"c0", (16384 + 856) => x"00", (16384 + 857) => x"ee", (16384 + 858) => x"71", (16384 + 859) => x"01", (16384 + 860) => x"13", (16384 + 861) => x"50", (16384 + 862) => x"60", (16384 + 863) => x"1b", (16384 + 864) => x"6b", (16384 + 865) => x"00", (16384 + 866) => x"d0", (16384 + 867) => x"11", (16384 + 868) => x"3f", (16384 + 869) => x"00", (16384 + 870) => x"7b", (16384 + 871) => x"01", (16384 + 872) => x"d0", (16384 + 873) => x"11", (16384 + 874) => x"70", (16384 + 875) => x"01", (16384 + 876) => x"30", (16384 + 877) => x"25", (16384 + 878) => x"13", (16384 + 879) => x"62", (16384 + 880) => x"00", (16384 + 881) => x"ee", (16384 + 882) => x"60", (16384 + 883) => x"1b", (16384 + 884) => x"d0", (16384 + 885) => x"11", (16384 + 886) => x"70", (16384 + 887) => x"01", (16384 + 888) => x"30", (16384 + 889) => x"25", (16384 + 890) => x"13", (16384 + 891) => x"74", (16384 + 892) => x"8e", (16384 + 893) => x"10", (16384 + 894) => x"8d", (16384 + 895) => x"e0", (16384 + 896) => x"7e", (16384 + 897) => x"ff", (16384 + 898) => x"60", (16384 + 899) => x"1b", (16384 + 900) => x"6b", (16384 + 901) => x"00", (16384 + 902) => x"d0", (16384 + 903) => x"e1", (16384 + 904) => x"3f", (16384 + 905) => x"00", (16384 + 906) => x"13", (16384 + 907) => x"90", (16384 + 908) => x"d0", (16384 + 909) => x"e1", (16384 + 910) => x"13", (16384 + 911) => x"94", (16384 + 912) => x"d0", (16384 + 913) => x"d1", (16384 + 914) => x"7b", (16384 + 915) => x"01", (16384 + 916) => x"70", (16384 + 917) => x"01", (16384 + 918) => x"30", (16384 + 919) => x"25", (16384 + 920) => x"13", (16384 + 921) => x"86", (16384 + 922) => x"4b", (16384 + 923) => x"00", (16384 + 924) => x"13", (16384 + 925) => x"a6", (16384 + 926) => x"7d", (16384 + 927) => x"ff", (16384 + 928) => x"7e", (16384 + 929) => x"ff", (16384 + 930) => x"3d", (16384 + 931) => x"01", (16384 + 932) => x"13", (16384 + 933) => x"82", (16384 + 934) => x"23", (16384 + 935) => x"c0", (16384 + 936) => x"3f", (16384 + 937) => x"01", (16384 + 938) => x"23", (16384 + 939) => x"c0", (16384 + 940) => x"7a", (16384 + 941) => x"01", (16384 + 942) => x"23", (16384 + 943) => x"c0", (16384 + 944) => x"80", (16384 + 945) => x"a0", (16384 + 946) => x"6d", (16384 + 947) => x"07", (16384 + 948) => x"80", (16384 + 949) => x"d2", (16384 + 950) => x"40", (16384 + 951) => x"04", (16384 + 952) => x"75", (16384 + 953) => x"fe", (16384 + 954) => x"45", (16384 + 955) => x"02", (16384 + 956) => x"65", (16384 + 957) => x"04", (16384 + 958) => x"00", (16384 + 959) => x"ee", (16384 + 960) => x"a7", (16384 + 961) => x"00", (16384 + 962) => x"f2", (16384 + 963) => x"55", (16384 + 964) => x"a8", (16384 + 965) => x"04", (16384 + 966) => x"fa", (16384 + 967) => x"33", (16384 + 968) => x"f2", (16384 + 969) => x"65", (16384 + 970) => x"f0", (16384 + 971) => x"29", (16384 + 972) => x"6d", (16384 + 973) => x"32", (16384 + 974) => x"6e", (16384 + 975) => x"00", (16384 + 976) => x"dd", (16384 + 977) => x"e5", (16384 + 978) => x"7d", (16384 + 979) => x"05", (16384 + 980) => x"f1", (16384 + 981) => x"29", (16384 + 982) => x"dd", (16384 + 983) => x"e5", (16384 + 984) => x"7d", (16384 + 985) => x"05", (16384 + 986) => x"f2", (16384 + 987) => x"29", (16384 + 988) => x"dd", (16384 + 989) => x"e5", (16384 + 990) => x"a7", (16384 + 991) => x"00", (16384 + 992) => x"f2", (16384 + 993) => x"65", (16384 + 994) => x"a2", (16384 + 995) => x"b4", (16384 + 996) => x"00", (16384 + 997) => x"ee", (16384 + 998) => x"6a", (16384 + 999) => x"00", (16384 + 1000) => x"60", (16384 + 1001) => x"19", (16384 + 1002) => x"00", (16384 + 1003) => x"ee", (16384 + 1004) => x"37", (16384 + 1005) => x"23", 
                                
                                -- Blitz by David Winter
                                (20480 + 128) => x"00", (20480 + 129) => x"00", 
                                (20480 + 130) => x"0D", (20480 + 131) => x"00",
                                (20480 + 132) => x"00", (20480 + 133) => x"00",
                                (20480 + 134) => x"00", (20480 + 135) => x"00",
                                (20480 + 136) => x"00", (20480 + 137) => x"20", -- delay
                                (20480 + 138) => x"00",
                                (20480 + 512) => x"12", (20480 + 513) => x"17", (20480 + 514) => x"42", (20480 + 515) => x"4c", (20480 + 516) => x"49", (20480 + 517) => x"54", (20480 + 518) => x"5a", (20480 + 519) => x"20", (20480 + 520) => x"42", (20480 + 521) => x"79", (20480 + 522) => x"20", (20480 + 523) => x"44", (20480 + 524) => x"61", (20480 + 525) => x"76", (20480 + 526) => x"69", (20480 + 527) => x"64", (20480 + 528) => x"20", (20480 + 529) => x"57", (20480 + 530) => x"49", (20480 + 531) => x"4e", (20480 + 532) => x"54", (20480 + 533) => x"45", (20480 + 534) => x"52", (20480 + 535) => x"a3", (20480 + 536) => x"41", (20480 + 537) => x"60", (20480 + 538) => x"04", (20480 + 539) => x"61", (20480 + 540) => x"09", (20480 + 541) => x"62", (20480 + 542) => x"0e", (20480 + 543) => x"67", (20480 + 544) => x"04", (20480 + 545) => x"d0", (20480 + 546) => x"1e", (20480 + 547) => x"f2", (20480 + 548) => x"1e", (20480 + 549) => x"70", (20480 + 550) => x"0c", (20480 + 551) => x"30", (20480 + 552) => x"40", (20480 + 553) => x"12", (20480 + 554) => x"21", (20480 + 555) => x"f0", (20480 + 556) => x"0a", (20480 + 557) => x"00", (20480 + 558) => x"e0", (20480 + 559) => x"22", (20480 + 560) => x"d9", (20480 + 561) => x"f0", (20480 + 562) => x"0a", (20480 + 563) => x"00", (20480 + 564) => x"e0", (20480 + 565) => x"8e", (20480 + 566) => x"70", (20480 + 567) => x"a3", (20480 + 568) => x"1e", (20480 + 569) => x"6b", (20480 + 570) => x"1f", (20480 + 571) => x"cc", (20480 + 572) => x"1f", (20480 + 573) => x"8c", (20480 + 574) => x"c4", (20480 + 575) => x"dc", (20480 + 576) => x"b2", (20480 + 577) => x"3f", (20480 + 578) => x"01", (20480 + 579) => x"12", (20480 + 580) => x"49", (20480 + 581) => x"dc", (20480 + 582) => x"b2", (20480 + 583) => x"12", (20480 + 584) => x"39", (20480 + 585) => x"ca", (20480 + 586) => x"07", (20480 + 587) => x"7a", (20480 + 588) => x"01", (20480 + 589) => x"7b", (20480 + 590) => x"fe", (20480 + 591) => x"dc", (20480 + 592) => x"b2", (20480 + 593) => x"7a", (20480 + 594) => x"ff", (20480 + 595) => x"3a", (20480 + 596) => x"00", (20480 + 597) => x"12", (20480 + 598) => x"4d", (20480 + 599) => x"7e", (20480 + 600) => x"ff", (20480 + 601) => x"3e", (20480 + 602) => x"00", (20480 + 603) => x"12", (20480 + 604) => x"39", (20480 + 605) => x"6b", (20480 + 606) => x"00", (20480 + 607) => x"8c", (20480 + 608) => x"70", (20480 + 609) => x"6d", (20480 + 610) => x"00", (20480 + 611) => x"6e", (20480 + 612) => x"00", (20480 + 613) => x"a3", (20480 + 614) => x"1b", (20480 + 615) => x"dd", (20480 + 616) => x"e3", (20480 + 617) => x"3f", (20480 + 618) => x"00", (20480 + 619) => x"12", (20480 + 620) => x"c1", (20480 + 621) => x"3b", (20480 + 622) => x"00", (20480 + 623) => x"12", (20480 + 624) => x"81", (20480 + 625) => x"60", (20480 + 626) => x"05", (20480 + 627) => x"e0", (20480 + 628) => x"9e", (20480 + 629) => x"12", (20480 + 630) => x"87", (20480 + 631) => x"6b", (20480 + 632) => x"01", (20480 + 633) => x"88", (20480 + 634) => x"d0", (20480 + 635) => x"78", (20480 + 636) => x"02", (20480 + 637) => x"89", (20480 + 638) => x"e0", (20480 + 639) => x"79", (20480 + 640) => x"03", (20480 + 641) => x"a3", (20480 + 642) => x"1e", (20480 + 643) => x"d8", (20480 + 644) => x"91", (20480 + 645) => x"81", (20480 + 646) => x"f0", (20480 + 647) => x"60", (20480 + 648) => x"05", (20480 + 649) => x"f0", (20480 + 650) => x"15", (20480 + 651) => x"f0", (20480 + 652) => x"07", (20480 + 653) => x"30", (20480 + 654) => x"00", (20480 + 655) => x"12", (20480 + 656) => x"8b", (20480 + 657) => x"3b", (20480 + 658) => x"01", (20480 + 659) => x"12", (20480 + 660) => x"ab", (20480 + 661) => x"a3", (20480 + 662) => x"1e", (20480 + 663) => x"31", (20480 + 664) => x"01", (20480 + 665) => x"d8", (20480 + 666) => x"91", (20480 + 667) => x"79", (20480 + 668) => x"01", (20480 + 669) => x"39", (20480 + 670) => x"20", (20480 + 671) => x"12", (20480 + 672) => x"ab", (20480 + 673) => x"6b", (20480 + 674) => x"00", (20480 + 675) => x"31", (20480 + 676) => x"00", (20480 + 677) => x"7c", (20480 + 678) => x"ff", (20480 + 679) => x"4c", (20480 + 680) => x"00", (20480 + 681) => x"12", (20480 + 682) => x"bb", (20480 + 683) => x"a3", (20480 + 684) => x"1b", (20480 + 685) => x"dd", (20480 + 686) => x"e3", (20480 + 687) => x"7d", (20480 + 688) => x"02", (20480 + 689) => x"3d", (20480 + 690) => x"40", (20480 + 691) => x"12", (20480 + 692) => x"b9", (20480 + 693) => x"6d", (20480 + 694) => x"00", (20480 + 695) => x"7e", (20480 + 696) => x"01", (20480 + 697) => x"12", (20480 + 698) => x"65", (20480 + 699) => x"00", (20480 + 700) => x"e0", (20480 + 701) => x"77", (20480 + 702) => x"02", (20480 + 703) => x"12", (20480 + 704) => x"2d", (20480 + 705) => x"a3", (20480 + 706) => x"1b", (20480 + 707) => x"dd", (20480 + 708) => x"e3", (20480 + 709) => x"60", (20480 + 710) => x"14", (20480 + 711) => x"61", (20480 + 712) => x"02", (20480 + 713) => x"62", (20480 + 714) => x"0b", (20480 + 715) => x"a3", (20480 + 716) => x"20", (20480 + 717) => x"d0", (20480 + 718) => x"1b", (20480 + 719) => x"f2", (20480 + 720) => x"1e", (20480 + 721) => x"70", (20480 + 722) => x"08", (20480 + 723) => x"30", (20480 + 724) => x"2c", (20480 + 725) => x"12", (20480 + 726) => x"cd", (20480 + 727) => x"12", (20480 + 728) => x"d7", (20480 + 729) => x"60", (20480 + 730) => x"0a", (20480 + 731) => x"61", (20480 + 732) => x"0d", (20480 + 733) => x"62", (20480 + 734) => x"05", (20480 + 735) => x"a3", (20480 + 736) => x"07", (20480 + 737) => x"d0", (20480 + 738) => x"15", (20480 + 739) => x"f2", (20480 + 740) => x"1e", (20480 + 741) => x"70", (20480 + 742) => x"08", (20480 + 743) => x"30", (20480 + 744) => x"2a", (20480 + 745) => x"12", (20480 + 746) => x"e1", (20480 + 747) => x"80", (20480 + 748) => x"70", (20480 + 749) => x"70", (20480 + 750) => x"fe", (20480 + 751) => x"80", (20480 + 752) => x"06", (20480 + 753) => x"a3", (20480 + 754) => x"87", (20480 + 755) => x"f0", (20480 + 756) => x"33", (20480 + 757) => x"f2", (20480 + 758) => x"65", (20480 + 759) => x"60", (20480 + 760) => x"2d", (20480 + 761) => x"f1", (20480 + 762) => x"29", (20480 + 763) => x"61", (20480 + 764) => x"0d", (20480 + 765) => x"d0", (20480 + 766) => x"15", (20480 + 767) => x"70", (20480 + 768) => x"05", (20480 + 769) => x"f2", (20480 + 770) => x"29", (20480 + 771) => x"d0", (20480 + 772) => x"15", (20480 + 773) => x"00", (20480 + 774) => x"ee", (20480 + 775) => x"83", (20480 + 776) => x"82", (20480 + 777) => x"83", (20480 + 778) => x"82", (20480 + 779) => x"fb", (20480 + 780) => x"e8", (20480 + 781) => x"08", (20480 + 782) => x"88", (20480 + 783) => x"05", (20480 + 784) => x"e2", (20480 + 785) => x"be", (20480 + 786) => x"a0", (20480 + 787) => x"b8", (20480 + 788) => x"20", (20480 + 789) => x"3e", (20480 + 790) => x"80", (20480 + 791) => x"80", (20480 + 792) => x"80", (20480 + 793) => x"80", (20480 + 794) => x"f8", (20480 + 795) => x"80", (20480 + 796) => x"f8", (20480 + 797) => x"fc", (20480 + 798) => x"c0", (20480 + 799) => x"c0", (20480 + 800) => x"f9", (20480 + 801) => x"81", (20480 + 802) => x"db", (20480 + 803) => x"cb", (20480 + 804) => x"fb", (20480 + 805) => x"00", (20480 + 806) => x"fa", (20480 + 807) => x"8a", (20480 + 808) => x"9a", (20480 + 809) => x"99", (20480 + 810) => x"f8", (20480 + 811) => x"ef", (20480 + 812) => x"2a", (20480 + 813) => x"e8", (20480 + 814) => x"29", (20480 + 815) => x"29", (20480 + 816) => x"00", (20480 + 817) => x"6f", (20480 + 818) => x"68", (20480 + 819) => x"2e", (20480 + 820) => x"4c", (20480 + 821) => x"8f", (20480 + 822) => x"be", (20480 + 823) => x"a0", (20480 + 824) => x"b8", (20480 + 825) => x"b0", (20480 + 826) => x"be", (20480 + 827) => x"00", (20480 + 828) => x"be", (20480 + 829) => x"22", (20480 + 830) => x"3e", (20480 + 831) => x"34", (20480 + 832) => x"b2", (20480 + 833) => x"d8", (20480 + 834) => x"d8", (20480 + 835) => x"00", (20480 + 836) => x"c3", (20480 + 837) => x"c3", (20480 + 838) => x"00", (20480 + 839) => x"d8", (20480 + 840) => x"d8", (20480 + 841) => x"00", (20480 + 842) => x"c3", (20480 + 843) => x"c3", (20480 + 844) => x"00", (20480 + 845) => x"d8", (20480 + 846) => x"d8", (20480 + 847) => x"c0", (20480 + 848) => x"c0", (20480 + 849) => x"00", (20480 + 850) => x"c0", (20480 + 851) => x"c0", (20480 + 852) => x"00", (20480 + 853) => x"c0", (20480 + 854) => x"c0", (20480 + 855) => x"00", (20480 + 856) => x"c0", (20480 + 857) => x"c0", (20480 + 858) => x"00", (20480 + 859) => x"db", (20480 + 860) => x"db", (20480 + 861) => x"db", (20480 + 862) => x"db", (20480 + 863) => x"00", (20480 + 864) => x"18", (20480 + 865) => x"18", (20480 + 866) => x"00", (20480 + 867) => x"18", (20480 + 868) => x"18", (20480 + 869) => x"00", (20480 + 870) => x"18", (20480 + 871) => x"18", (20480 + 872) => x"00", (20480 + 873) => x"db", (20480 + 874) => x"db", (20480 + 875) => x"db", (20480 + 876) => x"db", (20480 + 877) => x"00", (20480 + 878) => x"18", (20480 + 879) => x"18", (20480 + 880) => x"00", (20480 + 881) => x"18", (20480 + 882) => x"18", (20480 + 883) => x"00", (20480 + 884) => x"18", (20480 + 885) => x"18", (20480 + 886) => x"00", (20480 + 887) => x"18", (20480 + 888) => x"18", (20480 + 889) => x"db", (20480 + 890) => x"db", (20480 + 891) => x"00", (20480 + 892) => x"03", (20480 + 893) => x"03", (20480 + 894) => x"00", (20480 + 895) => x"18", (20480 + 896) => x"18", (20480 + 897) => x"00", (20480 + 898) => x"c0", (20480 + 899) => x"c0", (20480 + 900) => x"00", (20480 + 901) => x"db", (20480 + 902) => x"db", (20480 + 903) => x"00", 
                                
                                -- Brix by Andre Gustafsson
                                (24576 + 128) => x"00", (24576 + 129) => x"00", 
                                (24576 + 130) => x"C0", (24576 + 131) => x"E0",
                                (24576 + 132) => x"00", (24576 + 133) => x"00",
                                (24576 + 134) => x"00", (24576 + 135) => x"00",
                                (24576 + 136) => x"00", (24576 + 137) => x"30", -- delay
                                (24576 + 138) => x"00",
                                (24576 + 512) => x"6e", (24576 + 513) => x"05", (24576 + 514) => x"65", (24576 + 515) => x"00", (24576 + 516) => x"6b", (24576 + 517) => x"06", (24576 + 518) => x"6a", (24576 + 519) => x"00", (24576 + 520) => x"a3", (24576 + 521) => x"0c", (24576 + 522) => x"da", (24576 + 523) => x"b1", (24576 + 524) => x"7a", (24576 + 525) => x"04", (24576 + 526) => x"3a", (24576 + 527) => x"40", (24576 + 528) => x"12", (24576 + 529) => x"08", (24576 + 530) => x"7b", (24576 + 531) => x"02", (24576 + 532) => x"3b", (24576 + 533) => x"12", (24576 + 534) => x"12", (24576 + 535) => x"06", (24576 + 536) => x"6c", (24576 + 537) => x"20", (24576 + 538) => x"6d", (24576 + 539) => x"1f", (24576 + 540) => x"a3", (24576 + 541) => x"10", (24576 + 542) => x"dc", (24576 + 543) => x"d1", (24576 + 544) => x"22", (24576 + 545) => x"f6", (24576 + 546) => x"60", (24576 + 547) => x"00", (24576 + 548) => x"61", (24576 + 549) => x"00", (24576 + 550) => x"a3", (24576 + 551) => x"12", (24576 + 552) => x"d0", (24576 + 553) => x"11", (24576 + 554) => x"70", (24576 + 555) => x"08", (24576 + 556) => x"a3", (24576 + 557) => x"0e", (24576 + 558) => x"d0", (24576 + 559) => x"11", (24576 + 560) => x"60", (24576 + 561) => x"40", (24576 + 562) => x"f0", (24576 + 563) => x"15", (24576 + 564) => x"f0", (24576 + 565) => x"07", (24576 + 566) => x"30", (24576 + 567) => x"00", (24576 + 568) => x"12", (24576 + 569) => x"34", (24576 + 570) => x"c6", (24576 + 571) => x"0f", (24576 + 572) => x"67", (24576 + 573) => x"1e", (24576 + 574) => x"68", (24576 + 575) => x"01", (24576 + 576) => x"69", (24576 + 577) => x"ff", (24576 + 578) => x"a3", (24576 + 579) => x"0e", (24576 + 580) => x"d6", (24576 + 581) => x"71", (24576 + 582) => x"a3", (24576 + 583) => x"10", (24576 + 584) => x"dc", (24576 + 585) => x"d1", (24576 + 586) => x"60", (24576 + 587) => x"04", (24576 + 588) => x"e0", (24576 + 589) => x"a1", (24576 + 590) => x"7c", (24576 + 591) => x"fe", (24576 + 592) => x"60", (24576 + 593) => x"06", (24576 + 594) => x"e0", (24576 + 595) => x"a1", (24576 + 596) => x"7c", (24576 + 597) => x"02", (24576 + 598) => x"60", (24576 + 599) => x"3f", (24576 + 600) => x"8c", (24576 + 601) => x"02", (24576 + 602) => x"dc", (24576 + 603) => x"d1", (24576 + 604) => x"a3", (24576 + 605) => x"0e", (24576 + 606) => x"d6", (24576 + 607) => x"71", (24576 + 608) => x"86", (24576 + 609) => x"84", (24576 + 610) => x"87", (24576 + 611) => x"94", (24576 + 612) => x"60", (24576 + 613) => x"3f", (24576 + 614) => x"86", (24576 + 615) => x"02", (24576 + 616) => x"61", (24576 + 617) => x"1f", (24576 + 618) => x"87", (24576 + 619) => x"12", (24576 + 620) => x"47", (24576 + 621) => x"1f", (24576 + 622) => x"12", (24576 + 623) => x"ac", (24576 + 624) => x"46", (24576 + 625) => x"00", (24576 + 626) => x"68", (24576 + 627) => x"01", (24576 + 628) => x"46", (24576 + 629) => x"3f", (24576 + 630) => x"68", (24576 + 631) => x"ff", (24576 + 632) => x"47", (24576 + 633) => x"00", (24576 + 634) => x"69", (24576 + 635) => x"01", (24576 + 636) => x"d6", (24576 + 637) => x"71", (24576 + 638) => x"3f", (24576 + 639) => x"01", (24576 + 640) => x"12", (24576 + 641) => x"aa", (24576 + 642) => x"47", (24576 + 643) => x"1f", (24576 + 644) => x"12", (24576 + 645) => x"aa", (24576 + 646) => x"60", (24576 + 647) => x"05", (24576 + 648) => x"80", (24576 + 649) => x"75", (24576 + 650) => x"3f", (24576 + 651) => x"00", (24576 + 652) => x"12", (24576 + 653) => x"aa", (24576 + 654) => x"60", (24576 + 655) => x"01", (24576 + 656) => x"f0", (24576 + 657) => x"18", (24576 + 658) => x"80", (24576 + 659) => x"60", (24576 + 660) => x"61", (24576 + 661) => x"fc", (24576 + 662) => x"80", (24576 + 663) => x"12", (24576 + 664) => x"a3", (24576 + 665) => x"0c", (24576 + 666) => x"d0", (24576 + 667) => x"71", (24576 + 668) => x"60", (24576 + 669) => x"fe", (24576 + 670) => x"89", (24576 + 671) => x"03", (24576 + 672) => x"22", (24576 + 673) => x"f6", (24576 + 674) => x"75", (24576 + 675) => x"01", (24576 + 676) => x"22", (24576 + 677) => x"f6", (24576 + 678) => x"45", (24576 + 679) => x"60", (24576 + 680) => x"12", (24576 + 681) => x"de", (24576 + 682) => x"12", (24576 + 683) => x"46", (24576 + 684) => x"69", (24576 + 685) => x"ff", (24576 + 686) => x"80", (24576 + 687) => x"60", (24576 + 688) => x"80", (24576 + 689) => x"c5", (24576 + 690) => x"3f", (24576 + 691) => x"01", (24576 + 692) => x"12", (24576 + 693) => x"ca", (24576 + 694) => x"61", (24576 + 695) => x"02", (24576 + 696) => x"80", (24576 + 697) => x"15", (24576 + 698) => x"3f", (24576 + 699) => x"01", (24576 + 700) => x"12", (24576 + 701) => x"e0", (24576 + 702) => x"80", (24576 + 703) => x"15", (24576 + 704) => x"3f", (24576 + 705) => x"01", (24576 + 706) => x"12", (24576 + 707) => x"ee", (24576 + 708) => x"80", (24576 + 709) => x"15", (24576 + 710) => x"3f", (24576 + 711) => x"01", (24576 + 712) => x"12", (24576 + 713) => x"e8", (24576 + 714) => x"60", (24576 + 715) => x"20", (24576 + 716) => x"f0", (24576 + 717) => x"18", (24576 + 718) => x"a3", (24576 + 719) => x"0e", (24576 + 720) => x"7e", (24576 + 721) => x"ff", (24576 + 722) => x"80", (24576 + 723) => x"e0", (24576 + 724) => x"80", (24576 + 725) => x"04", (24576 + 726) => x"61", (24576 + 727) => x"00", (24576 + 728) => x"d0", (24576 + 729) => x"11", (24576 + 730) => x"3e", (24576 + 731) => x"00", (24576 + 732) => x"12", (24576 + 733) => x"30", (24576 + 734) => x"12", (24576 + 735) => x"de", (24576 + 736) => x"78", (24576 + 737) => x"ff", (24576 + 738) => x"48", (24576 + 739) => x"fe", (24576 + 740) => x"68", (24576 + 741) => x"ff", (24576 + 742) => x"12", (24576 + 743) => x"ee", (24576 + 744) => x"78", (24576 + 745) => x"01", (24576 + 746) => x"48", (24576 + 747) => x"02", (24576 + 748) => x"68", (24576 + 749) => x"01", (24576 + 750) => x"60", (24576 + 751) => x"04", (24576 + 752) => x"f0", (24576 + 753) => x"18", (24576 + 754) => x"69", (24576 + 755) => x"ff", (24576 + 756) => x"12", (24576 + 757) => x"70", (24576 + 758) => x"a3", (24576 + 759) => x"14", (24576 + 760) => x"f5", (24576 + 761) => x"33", (24576 + 762) => x"f2", (24576 + 763) => x"65", (24576 + 764) => x"f1", (24576 + 765) => x"29", (24576 + 766) => x"63", (24576 + 767) => x"37", (24576 + 768) => x"64", (24576 + 769) => x"00", (24576 + 770) => x"d3", (24576 + 771) => x"45", (24576 + 772) => x"73", (24576 + 773) => x"05", (24576 + 774) => x"f2", (24576 + 775) => x"29", (24576 + 776) => x"d3", (24576 + 777) => x"45", (24576 + 778) => x"00", (24576 + 779) => x"ee", (24576 + 780) => x"e0", (24576 + 781) => x"00", (24576 + 782) => x"80", (24576 + 783) => x"00", (24576 + 784) => x"fc", (24576 + 785) => x"00", (24576 + 786) => x"aa", (24576 + 787) => x"00", (24576 + 788) => x"00", (24576 + 789) => x"00", (24576 + 790) => x"00", (24576 + 791) => x"00", 
                                
                                -- Cave by 199x
                                (28672 + 128) => x"00", (28672 + 129) => x"B0", 
                                (28672 + 130) => x"C0", (28672 + 131) => x"E0",
                                (28672 + 132) => x"F0", (28672 + 133) => x"00",
                                (28672 + 134) => x"BE", (28672 + 135) => x"0D",
                                (28672 + 136) => x"00", (28672 + 137) => x"30", -- delay
                                (28672 + 138) => x"00",
                                (28672 + 512) => x"00", (28672 + 513) => x"e0", (28672 + 514) => x"64", (28672 + 515) => x"00", (28672 + 516) => x"65", (28672 + 517) => x"00", (28672 + 518) => x"a2", (28672 + 519) => x"0a", (28672 + 520) => x"12", (28672 + 521) => x"0c", (28672 + 522) => x"cc", (28672 + 523) => x"33", (28672 + 524) => x"66", (28672 + 525) => x"1e", (28672 + 526) => x"d4", (28672 + 527) => x"52", (28672 + 528) => x"d4", (28672 + 529) => x"62", (28672 + 530) => x"74", (28672 + 531) => x"08", (28672 + 532) => x"44", (28672 + 533) => x"40", (28672 + 534) => x"12", (28672 + 535) => x"1a", (28672 + 536) => x"12", (28672 + 537) => x"0e", (28672 + 538) => x"a2", (28672 + 539) => x"1e", (28672 + 540) => x"12", (28672 + 541) => x"2c", (28672 + 542) => x"ff", (28672 + 543) => x"ff", (28672 + 544) => x"c0", (28672 + 545) => x"c0", (28672 + 546) => x"c0", (28672 + 547) => x"c0", (28672 + 548) => x"c0", (28672 + 549) => x"c0", (28672 + 550) => x"c0", (28672 + 551) => x"c0", (28672 + 552) => x"c0", (28672 + 553) => x"c0", (28672 + 554) => x"ff", (28672 + 555) => x"ff", (28672 + 556) => x"64", (28672 + 557) => x"0d", (28672 + 558) => x"65", (28672 + 559) => x"09", (28672 + 560) => x"d4", (28672 + 561) => x"5e", (28672 + 562) => x"74", (28672 + 563) => x"0a", (28672 + 564) => x"a2", (28672 + 565) => x"3a", (28672 + 566) => x"d4", (28672 + 567) => x"5e", (28672 + 568) => x"12", (28672 + 569) => x"48", (28672 + 570) => x"ff", (28672 + 571) => x"ff", (28672 + 572) => x"c3", (28672 + 573) => x"c3", (28672 + 574) => x"c3", (28672 + 575) => x"c3", (28672 + 576) => x"c3", (28672 + 577) => x"ff", (28672 + 578) => x"ff", (28672 + 579) => x"c3", (28672 + 580) => x"c3", (28672 + 581) => x"c3", (28672 + 582) => x"c3", (28672 + 583) => x"c3", (28672 + 584) => x"74", (28672 + 585) => x"0a", (28672 + 586) => x"a2", (28672 + 587) => x"50", (28672 + 588) => x"d4", (28672 + 589) => x"5e", (28672 + 590) => x"12", (28672 + 591) => x"5e", (28672 + 592) => x"c3", (28672 + 593) => x"c3", (28672 + 594) => x"c3", (28672 + 595) => x"c3", (28672 + 596) => x"c3", (28672 + 597) => x"66", (28672 + 598) => x"66", (28672 + 599) => x"66", (28672 + 600) => x"66", (28672 + 601) => x"66", (28672 + 602) => x"3c", (28672 + 603) => x"3c", (28672 + 604) => x"18", (28672 + 605) => x"18", (28672 + 606) => x"74", (28672 + 607) => x"0a", (28672 + 608) => x"a2", (28672 + 609) => x"66", (28672 + 610) => x"d4", (28672 + 611) => x"5e", (28672 + 612) => x"12", (28672 + 613) => x"74", (28672 + 614) => x"ff", (28672 + 615) => x"ff", (28672 + 616) => x"c0", (28672 + 617) => x"c0", (28672 + 618) => x"c0", (28672 + 619) => x"c0", (28672 + 620) => x"ff", (28672 + 621) => x"ff", (28672 + 622) => x"c0", (28672 + 623) => x"c0", (28672 + 624) => x"c0", (28672 + 625) => x"c0", (28672 + 626) => x"ff", (28672 + 627) => x"ff", (28672 + 628) => x"6a", (28672 + 629) => x"01", (28672 + 630) => x"6b", (28672 + 631) => x"04", (28672 + 632) => x"6c", (28672 + 633) => x"0e", (28672 + 634) => x"6d", (28672 + 635) => x"00", (28672 + 636) => x"a2", (28672 + 637) => x"81", (28672 + 638) => x"12", (28672 + 639) => x"a6", (28672 + 640) => x"80", (28672 + 641) => x"ff", (28672 + 642) => x"ff", (28672 + 643) => x"ff", (28672 + 644) => x"ff", (28672 + 645) => x"ff", (28672 + 646) => x"ff", (28672 + 647) => x"ff", (28672 + 648) => x"ff", (28672 + 649) => x"ff", (28672 + 650) => x"00", (28672 + 651) => x"e0", (28672 + 652) => x"64", (28672 + 653) => x"00", (28672 + 654) => x"65", (28672 + 655) => x"00", (28672 + 656) => x"d4", (28672 + 657) => x"58", (28672 + 658) => x"74", (28672 + 659) => x"08", (28672 + 660) => x"44", (28672 + 661) => x"40", (28672 + 662) => x"22", (28672 + 663) => x"9e", (28672 + 664) => x"45", (28672 + 665) => x"20", (28672 + 666) => x"12", (28672 + 667) => x"a4", (28672 + 668) => x"12", (28672 + 669) => x"90", (28672 + 670) => x"64", (28672 + 671) => x"00", (28672 + 672) => x"75", (28672 + 673) => x"08", (28672 + 674) => x"00", (28672 + 675) => x"ee", (28672 + 676) => x"12", (28672 + 677) => x"ae", (28672 + 678) => x"60", (28672 + 679) => x"0f", (28672 + 680) => x"e0", (28672 + 681) => x"9e", (28672 + 682) => x"12", (28672 + 683) => x"a8", (28672 + 684) => x"12", (28672 + 685) => x"8a", (28672 + 686) => x"4a", (28672 + 687) => x"01", (28672 + 688) => x"22", (28672 + 689) => x"d0", (28672 + 690) => x"4a", (28672 + 691) => x"02", (28672 + 692) => x"23", (28672 + 693) => x"8a", (28672 + 694) => x"4a", (28672 + 695) => x"03", (28672 + 696) => x"23", (28672 + 697) => x"b8", (28672 + 698) => x"4a", (28672 + 699) => x"04", (28672 + 700) => x"23", (28672 + 701) => x"e0", (28672 + 702) => x"4a", (28672 + 703) => x"05", (28672 + 704) => x"24", (28672 + 705) => x"18", (28672 + 706) => x"4a", (28672 + 707) => x"06", (28672 + 708) => x"24", (28672 + 709) => x"78", (28672 + 710) => x"4a", (28672 + 711) => x"07", (28672 + 712) => x"24", (28672 + 713) => x"e6", (28672 + 714) => x"4a", (28672 + 715) => x"08", (28672 + 716) => x"25", (28672 + 717) => x"10", (28672 + 718) => x"13", (28672 + 719) => x"18", (28672 + 720) => x"a2", (28672 + 721) => x"81", (28672 + 722) => x"64", (28672 + 723) => x"02", (28672 + 724) => x"65", (28672 + 725) => x"02", (28672 + 726) => x"d4", (28672 + 727) => x"58", (28672 + 728) => x"65", (28672 + 729) => x"0a", (28672 + 730) => x"d4", (28672 + 731) => x"58", (28672 + 732) => x"65", (28672 + 733) => x"12", (28672 + 734) => x"d4", (28672 + 735) => x"58", (28672 + 736) => x"64", (28672 + 737) => x"0a", (28672 + 738) => x"65", (28672 + 739) => x"05", (28672 + 740) => x"d4", (28672 + 741) => x"53", (28672 + 742) => x"64", (28672 + 743) => x"12", (28672 + 744) => x"d4", (28672 + 745) => x"53", (28672 + 746) => x"64", (28672 + 747) => x"1a", (28672 + 748) => x"d4", (28672 + 749) => x"53", (28672 + 750) => x"64", (28672 + 751) => x"22", (28672 + 752) => x"d4", (28672 + 753) => x"53", (28672 + 754) => x"64", (28672 + 755) => x"2a", (28672 + 756) => x"d4", (28672 + 757) => x"53", (28672 + 758) => x"64", (28672 + 759) => x"32", (28672 + 760) => x"d4", (28672 + 761) => x"53", (28672 + 762) => x"a2", (28672 + 763) => x"fe", (28672 + 764) => x"13", (28672 + 765) => x"0a", (28672 + 766) => x"fc", (28672 + 767) => x"fc", (28672 + 768) => x"fc", (28672 + 769) => x"fc", (28672 + 770) => x"fc", (28672 + 771) => x"fc", (28672 + 772) => x"fc", (28672 + 773) => x"fc", (28672 + 774) => x"fc", (28672 + 775) => x"fc", (28672 + 776) => x"fc", (28672 + 777) => x"fc", (28672 + 778) => x"75", (28672 + 779) => x"03", (28672 + 780) => x"74", (28672 + 781) => x"02", (28672 + 782) => x"d4", (28672 + 783) => x"5c", (28672 + 784) => x"74", (28672 + 785) => x"06", (28672 + 786) => x"75", (28672 + 787) => x"09", (28672 + 788) => x"d4", (28672 + 789) => x"53", (28672 + 790) => x"00", (28672 + 791) => x"ee", (28672 + 792) => x"a2", (28672 + 793) => x"80", (28672 + 794) => x"db", (28672 + 795) => x"c1", (28672 + 796) => x"4f", (28672 + 797) => x"01", (28672 + 798) => x"13", (28672 + 799) => x"72", (28672 + 800) => x"60", (28672 + 801) => x"02", (28672 + 802) => x"e0", (28672 + 803) => x"a1", (28672 + 804) => x"6d", (28672 + 805) => x"02", (28672 + 806) => x"60", (28672 + 807) => x"04", (28672 + 808) => x"e0", (28672 + 809) => x"a1", (28672 + 810) => x"6d", (28672 + 811) => x"04", (28672 + 812) => x"60", (28672 + 813) => x"06", (28672 + 814) => x"e0", (28672 + 815) => x"a1", (28672 + 816) => x"6d", (28672 + 817) => x"06", (28672 + 818) => x"60", (28672 + 819) => x"08", (28672 + 820) => x"e0", (28672 + 821) => x"a1", (28672 + 822) => x"6d", (28672 + 823) => x"08", (28672 + 824) => x"db", (28672 + 825) => x"c1", (28672 + 826) => x"4d", (28672 + 827) => x"02", (28672 + 828) => x"7c", (28672 + 829) => x"ff", (28672 + 830) => x"4d", (28672 + 831) => x"04", (28672 + 832) => x"7b", (28672 + 833) => x"ff", (28672 + 834) => x"4d", (28672 + 835) => x"06", (28672 + 836) => x"7b", (28672 + 837) => x"01", (28672 + 838) => x"4d", (28672 + 839) => x"08", (28672 + 840) => x"7c", (28672 + 841) => x"01", (28672 + 842) => x"4b", (28672 + 843) => x"40", (28672 + 844) => x"13", (28672 + 845) => x"5e", (28672 + 846) => x"4b", (28672 + 847) => x"ff", (28672 + 848) => x"13", (28672 + 849) => x"64", (28672 + 850) => x"60", (28672 + 851) => x"02", (28672 + 852) => x"f0", (28672 + 853) => x"15", (28672 + 854) => x"f0", (28672 + 855) => x"07", (28672 + 856) => x"30", (28672 + 857) => x"00", (28672 + 858) => x"13", (28672 + 859) => x"56", (28672 + 860) => x"13", (28672 + 861) => x"18", (28672 + 862) => x"7a", (28672 + 863) => x"01", (28672 + 864) => x"4a", (28672 + 865) => x"09", (28672 + 866) => x"15", (28672 + 867) => x"3a", (28672 + 868) => x"6b", (28672 + 869) => x"01", (28672 + 870) => x"a2", (28672 + 871) => x"81", (28672 + 872) => x"12", (28672 + 873) => x"8a", (28672 + 874) => x"7a", (28672 + 875) => x"ff", (28672 + 876) => x"6b", (28672 + 877) => x"3e", (28672 + 878) => x"a2", (28672 + 879) => x"81", (28672 + 880) => x"12", (28672 + 881) => x"8a", (28672 + 882) => x"60", (28672 + 883) => x"03", (28672 + 884) => x"f0", (28672 + 885) => x"18", (28672 + 886) => x"60", (28672 + 887) => x"0f", (28672 + 888) => x"e0", (28672 + 889) => x"9e", (28672 + 890) => x"13", (28672 + 891) => x"78", (28672 + 892) => x"6a", (28672 + 893) => x"01", (28672 + 894) => x"6b", (28672 + 895) => x"04", (28672 + 896) => x"6c", (28672 + 897) => x"0e", (28672 + 898) => x"6d", (28672 + 899) => x"00", (28672 + 900) => x"a2", (28672 + 901) => x"81", (28672 + 902) => x"00", (28672 + 903) => x"e0", (28672 + 904) => x"12", (28672 + 905) => x"8a", (28672 + 906) => x"64", (28672 + 907) => x"00", (28672 + 908) => x"65", (28672 + 909) => x"11", (28672 + 910) => x"a2", (28672 + 911) => x"81", (28672 + 912) => x"d4", (28672 + 913) => x"53", (28672 + 914) => x"74", (28672 + 915) => x"08", (28672 + 916) => x"d4", (28672 + 917) => x"53", (28672 + 918) => x"74", (28672 + 919) => x"08", (28672 + 920) => x"75", (28672 + 921) => x"ff", (28672 + 922) => x"d4", (28672 + 923) => x"53", (28672 + 924) => x"74", (28672 + 925) => x"08", (28672 + 926) => x"75", (28672 + 927) => x"ff", (28672 + 928) => x"d4", (28672 + 929) => x"53", (28672 + 930) => x"74", (28672 + 931) => x"08", (28672 + 932) => x"d4", (28672 + 933) => x"53", (28672 + 934) => x"74", (28672 + 935) => x"08", (28672 + 936) => x"d4", (28672 + 937) => x"53", (28672 + 938) => x"74", (28672 + 939) => x"08", (28672 + 940) => x"75", (28672 + 941) => x"01", (28672 + 942) => x"d4", (28672 + 943) => x"53", (28672 + 944) => x"74", (28672 + 945) => x"08", (28672 + 946) => x"75", (28672 + 947) => x"01", (28672 + 948) => x"d4", (28672 + 949) => x"53", (28672 + 950) => x"00", (28672 + 951) => x"ee", (28672 + 952) => x"64", (28672 + 953) => x"00", (28672 + 954) => x"65", (28672 + 955) => x"11", (28672 + 956) => x"a2", (28672 + 957) => x"81", (28672 + 958) => x"d4", (28672 + 959) => x"53", (28672 + 960) => x"74", (28672 + 961) => x"08", (28672 + 962) => x"d4", (28672 + 963) => x"53", (28672 + 964) => x"74", (28672 + 965) => x"08", (28672 + 966) => x"75", (28672 + 967) => x"02", (28672 + 968) => x"d4", (28672 + 969) => x"52", (28672 + 970) => x"74", (28672 + 971) => x"08", (28672 + 972) => x"d4", (28672 + 973) => x"51", (28672 + 974) => x"74", (28672 + 975) => x"08", (28672 + 976) => x"d4", (28672 + 977) => x"51", (28672 + 978) => x"74", (28672 + 979) => x"08", (28672 + 980) => x"d4", (28672 + 981) => x"51", (28672 + 982) => x"74", (28672 + 983) => x"08", (28672 + 984) => x"d4", (28672 + 985) => x"51", (28672 + 986) => x"74", (28672 + 987) => x"08", (28672 + 988) => x"d4", (28672 + 989) => x"51", (28672 + 990) => x"00", (28672 + 991) => x"ee", (28672 + 992) => x"64", (28672 + 993) => x"00", (28672 + 994) => x"65", (28672 + 995) => x"13", (28672 + 996) => x"a2", (28672 + 997) => x"81", (28672 + 998) => x"d4", (28672 + 999) => x"51", (28672 + 1000) => x"a2", (28672 + 1001) => x"80", (28672 + 1002) => x"74", (28672 + 1003) => x"08", (28672 + 1004) => x"d4", (28672 + 1005) => x"51", (28672 + 1006) => x"75", (28672 + 1007) => x"01", (28672 + 1008) => x"d4", (28672 + 1009) => x"51", (28672 + 1010) => x"75", (28672 + 1011) => x"01", (28672 + 1012) => x"a2", (28672 + 1013) => x"81", (28672 + 1014) => x"d4", (28672 + 1015) => x"51", (28672 + 1016) => x"74", (28672 + 1017) => x"08", (28672 + 1018) => x"d4", (28672 + 1019) => x"51", (28672 + 1020) => x"74", (28672 + 1021) => x"08", (28672 + 1022) => x"d4", (28672 + 1023) => x"52", (28672 + 1024) => x"74", (28672 + 1025) => x"08", (28672 + 1026) => x"75", (28672 + 1027) => x"ff", (28672 + 1028) => x"d4", (28672 + 1029) => x"53", (28672 + 1030) => x"74", (28672 + 1031) => x"08", (28672 + 1032) => x"d4", (28672 + 1033) => x"54", (28672 + 1034) => x"74", (28672 + 1035) => x"08", (28672 + 1036) => x"75", (28672 + 1037) => x"ff", (28672 + 1038) => x"d4", (28672 + 1039) => x"56", (28672 + 1040) => x"74", (28672 + 1041) => x"08", (28672 + 1042) => x"75", (28672 + 1043) => x"ff", (28672 + 1044) => x"d4", (28672 + 1045) => x"58", (28672 + 1046) => x"00", (28672 + 1047) => x"ee", (28672 + 1048) => x"64", (28672 + 1049) => x"00", (28672 + 1050) => x"65", (28672 + 1051) => x"12", (28672 + 1052) => x"a2", (28672 + 1053) => x"81", (28672 + 1054) => x"d4", (28672 + 1055) => x"58", (28672 + 1056) => x"74", (28672 + 1057) => x"08", (28672 + 1058) => x"d4", (28672 + 1059) => x"58", (28672 + 1060) => x"74", (28672 + 1061) => x"08", (28672 + 1062) => x"d4", (28672 + 1063) => x"58", (28672 + 1064) => x"74", (28672 + 1065) => x"08", (28672 + 1066) => x"d4", (28672 + 1067) => x"58", (28672 + 1068) => x"74", (28672 + 1069) => x"08", (28672 + 1070) => x"d4", (28672 + 1071) => x"58", (28672 + 1072) => x"74", (28672 + 1073) => x"08", (28672 + 1074) => x"d4", (28672 + 1075) => x"58", (28672 + 1076) => x"74", (28672 + 1077) => x"08", (28672 + 1078) => x"d4", (28672 + 1079) => x"58", (28672 + 1080) => x"a2", (28672 + 1081) => x"80", (28672 + 1082) => x"75", (28672 + 1083) => x"ff", (28672 + 1084) => x"74", (28672 + 1085) => x"20", (28672 + 1086) => x"d4", (28672 + 1087) => x"51", (28672 + 1088) => x"75", (28672 + 1089) => x"ff", (28672 + 1090) => x"d4", (28672 + 1091) => x"51", (28672 + 1092) => x"75", (28672 + 1093) => x"ff", (28672 + 1094) => x"d4", (28672 + 1095) => x"51", (28672 + 1096) => x"75", (28672 + 1097) => x"ff", (28672 + 1098) => x"d4", (28672 + 1099) => x"51", (28672 + 1100) => x"75", (28672 + 1101) => x"ff", (28672 + 1102) => x"d4", (28672 + 1103) => x"51", (28672 + 1104) => x"75", (28672 + 1105) => x"ff", (28672 + 1106) => x"d4", (28672 + 1107) => x"51", (28672 + 1108) => x"75", (28672 + 1109) => x"ff", (28672 + 1110) => x"d4", (28672 + 1111) => x"51", (28672 + 1112) => x"75", (28672 + 1113) => x"ff", (28672 + 1114) => x"d4", (28672 + 1115) => x"51", (28672 + 1116) => x"75", (28672 + 1117) => x"ff", (28672 + 1118) => x"a2", (28672 + 1119) => x"81", (28672 + 1120) => x"d4", (28672 + 1121) => x"51", (28672 + 1122) => x"74", (28672 + 1123) => x"08", (28672 + 1124) => x"d4", (28672 + 1125) => x"51", (28672 + 1126) => x"74", (28672 + 1127) => x"08", (28672 + 1128) => x"d4", (28672 + 1129) => x"51", (28672 + 1130) => x"74", (28672 + 1131) => x"08", (28672 + 1132) => x"d4", (28672 + 1133) => x"51", (28672 + 1134) => x"74", (28672 + 1135) => x"08", (28672 + 1136) => x"d4", (28672 + 1137) => x"51", (28672 + 1138) => x"74", (28672 + 1139) => x"08", (28672 + 1140) => x"d4", (28672 + 1141) => x"51", (28672 + 1142) => x"00", (28672 + 1143) => x"ee", (28672 + 1144) => x"64", (28672 + 1145) => x"00", (28672 + 1146) => x"65", (28672 + 1147) => x"09", (28672 + 1148) => x"a2", (28672 + 1149) => x"81", (28672 + 1150) => x"d4", (28672 + 1151) => x"51", (28672 + 1152) => x"74", (28672 + 1153) => x"08", (28672 + 1154) => x"d4", (28672 + 1155) => x"51", (28672 + 1156) => x"74", (28672 + 1157) => x"08", (28672 + 1158) => x"d4", (28672 + 1159) => x"51", (28672 + 1160) => x"74", (28672 + 1161) => x"08", (28672 + 1162) => x"d4", (28672 + 1163) => x"51", (28672 + 1164) => x"74", (28672 + 1165) => x"08", (28672 + 1166) => x"d4", (28672 + 1167) => x"51", (28672 + 1168) => x"74", (28672 + 1169) => x"08", (28672 + 1170) => x"d4", (28672 + 1171) => x"51", (28672 + 1172) => x"a2", (28672 + 1173) => x"80", (28672 + 1174) => x"75", (28672 + 1175) => x"01", (28672 + 1176) => x"d4", (28672 + 1177) => x"51", (28672 + 1178) => x"75", (28672 + 1179) => x"01", (28672 + 1180) => x"d4", (28672 + 1181) => x"51", (28672 + 1182) => x"75", (28672 + 1183) => x"01", (28672 + 1184) => x"d4", (28672 + 1185) => x"51", (28672 + 1186) => x"75", (28672 + 1187) => x"01", (28672 + 1188) => x"d4", (28672 + 1189) => x"51", (28672 + 1190) => x"75", (28672 + 1191) => x"01", (28672 + 1192) => x"d4", (28672 + 1193) => x"51", (28672 + 1194) => x"75", (28672 + 1195) => x"01", (28672 + 1196) => x"d4", (28672 + 1197) => x"51", (28672 + 1198) => x"75", (28672 + 1199) => x"01", (28672 + 1200) => x"d4", (28672 + 1201) => x"51", (28672 + 1202) => x"75", (28672 + 1203) => x"01", (28672 + 1204) => x"d4", (28672 + 1205) => x"51", (28672 + 1206) => x"75", (28672 + 1207) => x"01", (28672 + 1208) => x"a2", (28672 + 1209) => x"81", (28672 + 1210) => x"d4", (28672 + 1211) => x"51", (28672 + 1212) => x"74", (28672 + 1213) => x"08", (28672 + 1214) => x"d4", (28672 + 1215) => x"51", (28672 + 1216) => x"74", (28672 + 1217) => x"08", (28672 + 1218) => x"d4", (28672 + 1219) => x"51", (28672 + 1220) => x"00", (28672 + 1221) => x"ee", (28672 + 1222) => x"64", (28672 + 1223) => x"00", (28672 + 1224) => x"65", (28672 + 1225) => x"1a", (28672 + 1226) => x"a2", (28672 + 1227) => x"81", (28672 + 1228) => x"d4", (28672 + 1229) => x"51", (28672 + 1230) => x"74", (28672 + 1231) => x"08", (28672 + 1232) => x"d4", (28672 + 1233) => x"51", (28672 + 1234) => x"74", (28672 + 1235) => x"08", (28672 + 1236) => x"d4", (28672 + 1237) => x"51", (28672 + 1238) => x"74", (28672 + 1239) => x"08", (28672 + 1240) => x"d4", (28672 + 1241) => x"51", (28672 + 1242) => x"74", (28672 + 1243) => x"08", (28672 + 1244) => x"d4", (28672 + 1245) => x"51", (28672 + 1246) => x"75", (28672 + 1247) => x"ff", (28672 + 1248) => x"d4", (28672 + 1249) => x"51", (28672 + 1250) => x"74", (28672 + 1251) => x"08", (28672 + 1252) => x"d4", (28672 + 1253) => x"51", (28672 + 1254) => x"74", (28672 + 1255) => x"08", (28672 + 1256) => x"d4", (28672 + 1257) => x"51", (28672 + 1258) => x"74", (28672 + 1259) => x"08", (28672 + 1260) => x"d4", (28672 + 1261) => x"51", (28672 + 1262) => x"00", (28672 + 1263) => x"ee", (28672 + 1264) => x"64", (28672 + 1265) => x"00", (28672 + 1266) => x"65", (28672 + 1267) => x"19", (28672 + 1268) => x"a2", (28672 + 1269) => x"81", (28672 + 1270) => x"d4", (28672 + 1271) => x"51", (28672 + 1272) => x"74", (28672 + 1273) => x"08", (28672 + 1274) => x"d4", (28672 + 1275) => x"51", (28672 + 1276) => x"74", (28672 + 1277) => x"08", (28672 + 1278) => x"d4", (28672 + 1279) => x"51", (28672 + 1280) => x"74", (28672 + 1281) => x"08", (28672 + 1282) => x"d4", (28672 + 1283) => x"51", (28672 + 1284) => x"74", (28672 + 1285) => x"08", (28672 + 1286) => x"d4", (28672 + 1287) => x"51", (28672 + 1288) => x"75", (28672 + 1289) => x"ff", (28672 + 1290) => x"d4", (28672 + 1291) => x"51", (28672 + 1292) => x"74", (28672 + 1293) => x"08", (28672 + 1294) => x"d4", (28672 + 1295) => x"51", (28672 + 1296) => x"74", (28672 + 1297) => x"08", (28672 + 1298) => x"d4", (28672 + 1299) => x"51", (28672 + 1300) => x"74", (28672 + 1301) => x"08", (28672 + 1302) => x"d4", (28672 + 1303) => x"51", (28672 + 1304) => x"00", (28672 + 1305) => x"ee", (28672 + 1306) => x"00", (28672 + 1307) => x"e0", (28672 + 1308) => x"67", (28672 + 1309) => x"03", (28672 + 1310) => x"68", (28672 + 1311) => x"03", (28672 + 1312) => x"a5", (28672 + 1313) => x"44", (28672 + 1314) => x"15", (28672 + 1315) => x"5c", (28672 + 1316) => x"ae", (28672 + 1317) => x"aa", (28672 + 1318) => x"ea", (28672 + 1319) => x"4a", (28672 + 1320) => x"4e", (28672 + 1321) => x"00", (28672 + 1322) => x"a4", (28672 + 1323) => x"a4", (28672 + 1324) => x"a4", (28672 + 1325) => x"a5", (28672 + 1326) => x"e2", (28672 + 1327) => x"00", (28672 + 1328) => x"5d", (28672 + 1329) => x"55", (28672 + 1330) => x"55", (28672 + 1331) => x"55", (28672 + 1332) => x"9d", (28672 + 1333) => x"00", (28672 + 1334) => x"c8", (28672 + 1335) => x"48", (28672 + 1336) => x"48", (28672 + 1337) => x"40", (28672 + 1338) => x"48", (28672 + 1339) => x"00", (28672 + 1340) => x"d7", (28672 + 1341) => x"85", (28672 + 1342) => x"a5", (28672 + 1343) => x"4a", (28672 + 1344) => x"77", (28672 + 1345) => x"08", (28672 + 1346) => x"d7", (28672 + 1347) => x"85", (28672 + 1348) => x"77", (28672 + 1349) => x"08", (28672 + 1350) => x"a5", (28672 + 1351) => x"50", (28672 + 1352) => x"d7", (28672 + 1353) => x"85", (28672 + 1354) => x"77", (28672 + 1355) => x"08", (28672 + 1356) => x"a5", (28672 + 1357) => x"56", (28672 + 1358) => x"d7", (28672 + 1359) => x"85", (28672 + 1360) => x"15", (28672 + 1361) => x"70", 
                                
                                -- Hidden by David Winter
                                (32768 + 128) => x"00", (32768 + 129) => x"B0", 
                                (32768 + 130) => x"CD", (32768 + 131) => x"E0",
                                (32768 + 132) => x"F0", (32768 + 133) => x"00",
                                (32768 + 134) => x"BE", (32768 + 135) => x"00",
                                (32768 + 136) => x"00", (32768 + 137) => x"60", -- delay
                                (32768 + 138) => x"00",
                                (32768 + 512) => x"12", (32768 + 513) => x"1d", (32768 + 514) => x"48", (32768 + 515) => x"49", (32768 + 516) => x"44", (32768 + 517) => x"44", (32768 + 518) => x"45", (32768 + 519) => x"4e", (32768 + 520) => x"21", (32768 + 521) => x"20", (32768 + 522) => x"31", (32768 + 523) => x"2e", (32768 + 524) => x"30", (32768 + 525) => x"20", (32768 + 526) => x"42", (32768 + 527) => x"79", (32768 + 528) => x"20", (32768 + 529) => x"44", (32768 + 530) => x"61", (32768 + 531) => x"76", (32768 + 532) => x"69", (32768 + 533) => x"64", (32768 + 534) => x"20", (32768 + 535) => x"57", (32768 + 536) => x"49", (32768 + 537) => x"4e", (32768 + 538) => x"54", (32768 + 539) => x"45", (32768 + 540) => x"52", (32768 + 541) => x"a4", (32768 + 542) => x"3f", (32768 + 543) => x"60", (32768 + 544) => x"00", (32768 + 545) => x"61", (32768 + 546) => x"40", (32768 + 547) => x"f1", (32768 + 548) => x"55", (32768 + 549) => x"a4", (32768 + 550) => x"3f", (32768 + 551) => x"60", (32768 + 552) => x"00", (32768 + 553) => x"f0", (32768 + 554) => x"55", (32768 + 555) => x"00", (32768 + 556) => x"e0", (32768 + 557) => x"a4", (32768 + 558) => x"7e", (32768 + 559) => x"60", (32768 + 560) => x"0c", (32768 + 561) => x"61", (32768 + 562) => x"08", (32768 + 563) => x"62", (32768 + 564) => x"0f", (32768 + 565) => x"d0", (32768 + 566) => x"1f", (32768 + 567) => x"70", (32768 + 568) => x"08", (32768 + 569) => x"f2", (32768 + 570) => x"1e", (32768 + 571) => x"30", (32768 + 572) => x"34", (32768 + 573) => x"12", (32768 + 574) => x"35", (32768 + 575) => x"f0", (32768 + 576) => x"0a", (32768 + 577) => x"00", (32768 + 578) => x"e0", (32768 + 579) => x"a4", (32768 + 580) => x"c9", (32768 + 581) => x"60", (32768 + 582) => x"13", (32768 + 583) => x"61", (32768 + 584) => x"0d", (32768 + 585) => x"62", (32768 + 586) => x"04", (32768 + 587) => x"d0", (32768 + 588) => x"14", (32768 + 589) => x"70", (32768 + 590) => x"08", (32768 + 591) => x"f2", (32768 + 592) => x"1e", (32768 + 593) => x"30", (32768 + 594) => x"2b", (32768 + 595) => x"12", (32768 + 596) => x"4b", (32768 + 597) => x"a4", (32768 + 598) => x"1f", (32768 + 599) => x"ff", (32768 + 600) => x"65", (32768 + 601) => x"a4", (32768 + 602) => x"2f", (32768 + 603) => x"ff", (32768 + 604) => x"55", (32768 + 605) => x"63", (32768 + 606) => x"40", (32768 + 607) => x"66", (32768 + 608) => x"08", (32768 + 609) => x"c1", (32768 + 610) => x"0f", (32768 + 611) => x"c2", (32768 + 612) => x"0f", (32768 + 613) => x"a4", (32768 + 614) => x"2f", (32768 + 615) => x"f1", (32768 + 616) => x"1e", (32768 + 617) => x"f0", (32768 + 618) => x"65", (32768 + 619) => x"84", (32768 + 620) => x"00", (32768 + 621) => x"a4", (32768 + 622) => x"2f", (32768 + 623) => x"f2", (32768 + 624) => x"1e", (32768 + 625) => x"f0", (32768 + 626) => x"65", (32768 + 627) => x"85", (32768 + 628) => x"00", (32768 + 629) => x"80", (32768 + 630) => x"40", (32768 + 631) => x"f0", (32768 + 632) => x"55", (32768 + 633) => x"a4", (32768 + 634) => x"2f", (32768 + 635) => x"f1", (32768 + 636) => x"1e", (32768 + 637) => x"80", (32768 + 638) => x"50", (32768 + 639) => x"f0", (32768 + 640) => x"55", (32768 + 641) => x"73", (32768 + 642) => x"ff", (32768 + 643) => x"33", (32768 + 644) => x"00", (32768 + 645) => x"12", (32768 + 646) => x"61", (32768 + 647) => x"00", (32768 + 648) => x"e0", (32768 + 649) => x"60", (32768 + 650) => x"00", (32768 + 651) => x"61", (32768 + 652) => x"00", (32768 + 653) => x"a4", (32768 + 654) => x"77", (32768 + 655) => x"d0", (32768 + 656) => x"17", (32768 + 657) => x"70", (32768 + 658) => x"08", (32768 + 659) => x"30", (32768 + 660) => x"20", (32768 + 661) => x"12", (32768 + 662) => x"8f", (32768 + 663) => x"60", (32768 + 664) => x"00", (32768 + 665) => x"71", (32768 + 666) => x"08", (32768 + 667) => x"31", (32768 + 668) => x"20", (32768 + 669) => x"12", (32768 + 670) => x"8f", (32768 + 671) => x"6c", (32768 + 672) => x"00", (32768 + 673) => x"6d", (32768 + 674) => x"00", (32768 + 675) => x"6e", (32768 + 676) => x"00", (32768 + 677) => x"a4", (32768 + 678) => x"3f", (32768 + 679) => x"f0", (32768 + 680) => x"65", (32768 + 681) => x"70", (32768 + 682) => x"01", (32768 + 683) => x"f0", (32768 + 684) => x"55", (32768 + 685) => x"23", (32768 + 686) => x"b9", (32768 + 687) => x"6a", (32768 + 688) => x"10", (32768 + 689) => x"23", (32768 + 690) => x"5d", (32768 + 691) => x"23", (32768 + 692) => x"cd", (32768 + 693) => x"8a", (32768 + 694) => x"90", (32768 + 695) => x"87", (32768 + 696) => x"d0", (32768 + 697) => x"88", (32768 + 698) => x"e0", (32768 + 699) => x"23", (32768 + 700) => x"5d", (32768 + 701) => x"23", (32768 + 702) => x"cd", (32768 + 703) => x"23", (32768 + 704) => x"b9", (32768 + 705) => x"a4", (32768 + 706) => x"2f", (32768 + 707) => x"f9", (32768 + 708) => x"1e", (32768 + 709) => x"f0", (32768 + 710) => x"65", (32768 + 711) => x"81", (32768 + 712) => x"00", (32768 + 713) => x"a4", (32768 + 714) => x"2f", (32768 + 715) => x"fa", (32768 + 716) => x"1e", (32768 + 717) => x"f0", (32768 + 718) => x"65", (32768 + 719) => x"50", (32768 + 720) => x"10", (32768 + 721) => x"13", (32768 + 722) => x"2b", (32768 + 723) => x"23", (32768 + 724) => x"df", (32768 + 725) => x"60", (32768 + 726) => x"20", (32768 + 727) => x"24", (32768 + 728) => x"01", (32768 + 729) => x"23", (32768 + 730) => x"df", (32768 + 731) => x"60", (32768 + 732) => x"00", (32768 + 733) => x"a4", (32768 + 734) => x"2f", (32768 + 735) => x"f9", (32768 + 736) => x"1e", (32768 + 737) => x"f0", (32768 + 738) => x"55", (32768 + 739) => x"a4", (32768 + 740) => x"2f", (32768 + 741) => x"fa", (32768 + 742) => x"1e", (32768 + 743) => x"f0", (32768 + 744) => x"55", (32768 + 745) => x"76", (32768 + 746) => x"ff", (32768 + 747) => x"36", (32768 + 748) => x"00", (32768 + 749) => x"12", (32768 + 750) => x"a5", (32768 + 751) => x"a4", (32768 + 752) => x"3f", (32768 + 753) => x"f1", (32768 + 754) => x"65", (32768 + 755) => x"82", (32768 + 756) => x"00", (32768 + 757) => x"80", (32768 + 758) => x"15", (32768 + 759) => x"3f", (32768 + 760) => x"00", (32768 + 761) => x"13", (32768 + 762) => x"01", (32768 + 763) => x"80", (32768 + 764) => x"20", (32768 + 765) => x"81", (32768 + 766) => x"20", (32768 + 767) => x"f1", (32768 + 768) => x"55", (32768 + 769) => x"00", (32768 + 770) => x"e0", (32768 + 771) => x"a5", (32768 + 772) => x"19", (32768 + 773) => x"60", (32768 + 774) => x"10", (32768 + 775) => x"61", (32768 + 776) => x"07", (32768 + 777) => x"62", (32768 + 778) => x"0e", (32768 + 779) => x"d0", (32768 + 780) => x"1f", (32768 + 781) => x"70", (32768 + 782) => x"08", (32768 + 783) => x"f2", (32768 + 784) => x"1e", (32768 + 785) => x"30", (32768 + 786) => x"30", (32768 + 787) => x"13", (32768 + 788) => x"0b", (32768 + 789) => x"a4", (32768 + 790) => x"3f", (32768 + 791) => x"f1", (32768 + 792) => x"65", (32768 + 793) => x"84", (32768 + 794) => x"10", (32768 + 795) => x"83", (32768 + 796) => x"00", (32768 + 797) => x"66", (32768 + 798) => x"09", (32768 + 799) => x"24", (32768 + 800) => x"0b", (32768 + 801) => x"66", (32768 + 802) => x"0f", (32768 + 803) => x"83", (32768 + 804) => x"40", (32768 + 805) => x"24", (32768 + 806) => x"0b", (32768 + 807) => x"f0", (32768 + 808) => x"0a", (32768 + 809) => x"12", (32768 + 810) => x"25", (32768 + 811) => x"23", (32768 + 812) => x"db", (32768 + 813) => x"60", (32768 + 814) => x"80", (32768 + 815) => x"24", (32768 + 816) => x"01", (32768 + 817) => x"23", (32768 + 818) => x"db", (32768 + 819) => x"a4", (32768 + 820) => x"2f", (32768 + 821) => x"fa", (32768 + 822) => x"1e", (32768 + 823) => x"f0", (32768 + 824) => x"65", (32768 + 825) => x"70", (32768 + 826) => x"ff", (32768 + 827) => x"23", (32768 + 828) => x"f3", (32768 + 829) => x"a4", (32768 + 830) => x"41", (32768 + 831) => x"f0", (32768 + 832) => x"1e", (32768 + 833) => x"d7", (32768 + 834) => x"87", (32768 + 835) => x"a4", (32768 + 836) => x"77", (32768 + 837) => x"d7", (32768 + 838) => x"87", (32768 + 839) => x"a4", (32768 + 840) => x"2f", (32768 + 841) => x"f9", (32768 + 842) => x"1e", (32768 + 843) => x"f0", (32768 + 844) => x"65", (32768 + 845) => x"70", (32768 + 846) => x"ff", (32768 + 847) => x"23", (32768 + 848) => x"f3", (32768 + 849) => x"a4", (32768 + 850) => x"41", (32768 + 851) => x"f0", (32768 + 852) => x"1e", (32768 + 853) => x"dd", (32768 + 854) => x"e7", (32768 + 855) => x"a4", (32768 + 856) => x"77", (32768 + 857) => x"dd", (32768 + 858) => x"e7", (32768 + 859) => x"12", (32768 + 860) => x"a5", (32768 + 861) => x"a4", (32768 + 862) => x"71", (32768 + 863) => x"dd", (32768 + 864) => x"e7", (32768 + 865) => x"fb", (32768 + 866) => x"0a", (32768 + 867) => x"dd", (32768 + 868) => x"e7", (32768 + 869) => x"3b", (32768 + 870) => x"04", (32768 + 871) => x"13", (32768 + 872) => x"71", (32768 + 873) => x"4d", (32768 + 874) => x"00", (32768 + 875) => x"13", (32768 + 876) => x"5d", (32768 + 877) => x"7d", (32768 + 878) => x"f8", (32768 + 879) => x"7c", (32768 + 880) => x"ff", (32768 + 881) => x"3b", (32768 + 882) => x"06", (32768 + 883) => x"13", (32768 + 884) => x"7d", (32768 + 885) => x"4d", (32768 + 886) => x"18", (32768 + 887) => x"13", (32768 + 888) => x"5d", (32768 + 889) => x"7d", (32768 + 890) => x"08", (32768 + 891) => x"7c", (32768 + 892) => x"01", (32768 + 893) => x"3b", (32768 + 894) => x"02", (32768 + 895) => x"13", (32768 + 896) => x"89", (32768 + 897) => x"4e", (32768 + 898) => x"00", (32768 + 899) => x"13", (32768 + 900) => x"5d", (32768 + 901) => x"7e", (32768 + 902) => x"f8", (32768 + 903) => x"7c", (32768 + 904) => x"fc", (32768 + 905) => x"3b", (32768 + 906) => x"08", (32768 + 907) => x"13", (32768 + 908) => x"95", (32768 + 909) => x"4e", (32768 + 910) => x"18", (32768 + 911) => x"13", (32768 + 912) => x"5d", (32768 + 913) => x"7e", (32768 + 914) => x"08", (32768 + 915) => x"7c", (32768 + 916) => x"04", (32768 + 917) => x"3b", (32768 + 918) => x"05", (32768 + 919) => x"13", (32768 + 920) => x"5d", (32768 + 921) => x"a4", (32768 + 922) => x"2f", (32768 + 923) => x"fc", (32768 + 924) => x"1e", (32768 + 925) => x"f0", (32768 + 926) => x"65", (32768 + 927) => x"40", (32768 + 928) => x"00", (32768 + 929) => x"13", (32768 + 930) => x"5d", (32768 + 931) => x"89", (32768 + 932) => x"c0", (32768 + 933) => x"99", (32768 + 934) => x"a0", (32768 + 935) => x"13", (32768 + 936) => x"5d", (32768 + 937) => x"70", (32768 + 938) => x"ff", (32768 + 939) => x"a4", (32768 + 940) => x"77", (32768 + 941) => x"dd", (32768 + 942) => x"e7", (32768 + 943) => x"a4", (32768 + 944) => x"41", (32768 + 945) => x"23", (32768 + 946) => x"f3", (32768 + 947) => x"f0", (32768 + 948) => x"1e", (32768 + 949) => x"dd", (32768 + 950) => x"e7", (32768 + 951) => x"00", (32768 + 952) => x"ee", (32768 + 953) => x"a4", (32768 + 954) => x"d5", (32768 + 955) => x"60", (32768 + 956) => x"24", (32768 + 957) => x"61", (32768 + 958) => x"0a", (32768 + 959) => x"62", (32768 + 960) => x"0b", (32768 + 961) => x"d0", (32768 + 962) => x"1b", (32768 + 963) => x"70", (32768 + 964) => x"08", (32768 + 965) => x"f2", (32768 + 966) => x"1e", (32768 + 967) => x"30", (32768 + 968) => x"3c", (32768 + 969) => x"13", (32768 + 970) => x"c1", (32768 + 971) => x"00", (32768 + 972) => x"ee", (32768 + 973) => x"60", (32768 + 974) => x"34", (32768 + 975) => x"61", (32768 + 976) => x"10", (32768 + 977) => x"a4", (32768 + 978) => x"f1", (32768 + 979) => x"d0", (32768 + 980) => x"15", (32768 + 981) => x"a4", (32768 + 982) => x"f6", (32768 + 983) => x"d0", (32768 + 984) => x"15", (32768 + 985) => x"00", (32768 + 986) => x"ee", (32768 + 987) => x"a4", (32768 + 988) => x"fb", (32768 + 989) => x"13", (32768 + 990) => x"e1", (32768 + 991) => x"a5", (32768 + 992) => x"0a", (32768 + 993) => x"60", (32768 + 994) => x"24", (32768 + 995) => x"61", (32768 + 996) => x"0d", (32768 + 997) => x"62", (32768 + 998) => x"05", (32768 + 999) => x"d0", (32768 + 1000) => x"15", (32768 + 1001) => x"70", (32768 + 1002) => x"08", (32768 + 1003) => x"f2", (32768 + 1004) => x"1e", (32768 + 1005) => x"30", (32768 + 1006) => x"3c", (32768 + 1007) => x"13", (32768 + 1008) => x"e7", (32768 + 1009) => x"00", (32768 + 1010) => x"ee", (32768 + 1011) => x"81", (32768 + 1012) => x"00", (32768 + 1013) => x"81", (32768 + 1014) => x"14", (32768 + 1015) => x"80", (32768 + 1016) => x"04", (32768 + 1017) => x"80", (32768 + 1018) => x"04", (32768 + 1019) => x"80", (32768 + 1020) => x"04", (32768 + 1021) => x"80", (32768 + 1022) => x"15", (32768 + 1023) => x"00", (32768 + 1024) => x"ee", (32768 + 1025) => x"f0", (32768 + 1026) => x"15", (32768 + 1027) => x"f0", (32768 + 1028) => x"07", (32768 + 1029) => x"30", (32768 + 1030) => x"00", (32768 + 1031) => x"14", (32768 + 1032) => x"03", (32768 + 1033) => x"00", (32768 + 1034) => x"ee", (32768 + 1035) => x"a4", (32768 + 1036) => x"2f", (32768 + 1037) => x"f3", (32768 + 1038) => x"33", (32768 + 1039) => x"f2", (32768 + 1040) => x"65", (32768 + 1041) => x"65", (32768 + 1042) => x"23", (32768 + 1043) => x"f1", (32768 + 1044) => x"29", (32768 + 1045) => x"d5", (32768 + 1046) => x"65", (32768 + 1047) => x"65", (32768 + 1048) => x"28", (32768 + 1049) => x"f2", (32768 + 1050) => x"29", (32768 + 1051) => x"d5", (32768 + 1052) => x"65", (32768 + 1053) => x"00", (32768 + 1054) => x"ee", (32768 + 1055) => x"01", (32768 + 1056) => x"02", (32768 + 1057) => x"03", (32768 + 1058) => x"04", (32768 + 1059) => x"08", (32768 + 1060) => x"07", (32768 + 1061) => x"06", (32768 + 1062) => x"05", (32768 + 1063) => x"05", (32768 + 1064) => x"06", (32768 + 1065) => x"07", (32768 + 1066) => x"08", (32768 + 1067) => x"04", (32768 + 1068) => x"03", (32768 + 1069) => x"02", (32768 + 1070) => x"01", (32768 + 1071) => x"01", (32768 + 1072) => x"02", (32768 + 1073) => x"03", (32768 + 1074) => x"04", (32768 + 1075) => x"08", (32768 + 1076) => x"07", (32768 + 1077) => x"06", (32768 + 1078) => x"05", (32768 + 1079) => x"05", (32768 + 1080) => x"06", (32768 + 1081) => x"07", (32768 + 1082) => x"08", (32768 + 1083) => x"04", (32768 + 1084) => x"03", (32768 + 1085) => x"02", (32768 + 1086) => x"01", (32768 + 1087) => x"00", (32768 + 1088) => x"00", (32768 + 1089) => x"fe", (32768 + 1090) => x"ee", (32768 + 1091) => x"c6", (32768 + 1092) => x"82", (32768 + 1093) => x"c6", (32768 + 1094) => x"ee", (32768 + 1095) => x"fe", (32768 + 1096) => x"fe", (32768 + 1097) => x"c6", (32768 + 1098) => x"c6", (32768 + 1099) => x"c6", (32768 + 1100) => x"fe", (32768 + 1101) => x"fe", (32768 + 1102) => x"c6", (32768 + 1103) => x"aa", (32768 + 1104) => x"82", (32768 + 1105) => x"aa", (32768 + 1106) => x"c6", (32768 + 1107) => x"fe", (32768 + 1108) => x"c6", (32768 + 1109) => x"82", (32768 + 1110) => x"82", (32768 + 1111) => x"82", (32768 + 1112) => x"c6", (32768 + 1113) => x"fe", (32768 + 1114) => x"ba", (32768 + 1115) => x"d6", (32768 + 1116) => x"ee", (32768 + 1117) => x"d6", (32768 + 1118) => x"ba", (32768 + 1119) => x"fe", (32768 + 1120) => x"ee", (32768 + 1121) => x"ee", (32768 + 1122) => x"82", (32768 + 1123) => x"ee", (32768 + 1124) => x"ee", (32768 + 1125) => x"fe", (32768 + 1126) => x"82", (32768 + 1127) => x"fe", (32768 + 1128) => x"82", (32768 + 1129) => x"fe", (32768 + 1130) => x"82", (32768 + 1131) => x"fe", (32768 + 1132) => x"aa", (32768 + 1133) => x"aa", (32768 + 1134) => x"aa", (32768 + 1135) => x"aa", (32768 + 1136) => x"aa", (32768 + 1137) => x"fe", (32768 + 1138) => x"fe", (32768 + 1139) => x"fe", (32768 + 1140) => x"fe", (32768 + 1141) => x"fe", (32768 + 1142) => x"fe", (32768 + 1143) => x"fe", (32768 + 1144) => x"aa", (32768 + 1145) => x"d6", (32768 + 1146) => x"aa", (32768 + 1147) => x"d6", (32768 + 1148) => x"aa", (32768 + 1149) => x"fe", (32768 + 1150) => x"8b", (32768 + 1151) => x"88", (32768 + 1152) => x"f8", (32768 + 1153) => x"88", (32768 + 1154) => x"8b", (32768 + 1155) => x"00", (32768 + 1156) => x"00", (32768 + 1157) => x"00", (32768 + 1158) => x"00", (32768 + 1159) => x"00", (32768 + 1160) => x"f0", (32768 + 1161) => x"48", (32768 + 1162) => x"48", (32768 + 1163) => x"48", (32768 + 1164) => x"f2", (32768 + 1165) => x"ef", (32768 + 1166) => x"84", (32768 + 1167) => x"84", (32768 + 1168) => x"84", (32768 + 1169) => x"ef", (32768 + 1170) => x"00", (32768 + 1171) => x"08", (32768 + 1172) => x"08", (32768 + 1173) => x"0a", (32768 + 1174) => x"00", (32768 + 1175) => x"8a", (32768 + 1176) => x"8a", (32768 + 1177) => x"aa", (32768 + 1178) => x"aa", (32768 + 1179) => x"52", (32768 + 1180) => x"3c", (32768 + 1181) => x"92", (32768 + 1182) => x"92", (32768 + 1183) => x"92", (32768 + 1184) => x"3c", (32768 + 1185) => x"00", (32768 + 1186) => x"e2", (32768 + 1187) => x"a3", (32768 + 1188) => x"e3", (32768 + 1189) => x"00", (32768 + 1190) => x"8b", (32768 + 1191) => x"c8", (32768 + 1192) => x"a8", (32768 + 1193) => x"98", (32768 + 1194) => x"88", (32768 + 1195) => x"fa", (32768 + 1196) => x"83", (32768 + 1197) => x"e2", (32768 + 1198) => x"82", (32768 + 1199) => x"fa", (32768 + 1200) => x"00", (32768 + 1201) => x"28", (32768 + 1202) => x"b8", (32768 + 1203) => x"90", (32768 + 1204) => x"00", (32768 + 1205) => x"ef", (32768 + 1206) => x"88", (32768 + 1207) => x"8e", (32768 + 1208) => x"88", (32768 + 1209) => x"8f", (32768 + 1210) => x"21", (32768 + 1211) => x"21", (32768 + 1212) => x"a1", (32768 + 1213) => x"60", (32768 + 1214) => x"21", (32768 + 1215) => x"00", (32768 + 1216) => x"00", (32768 + 1217) => x"00", (32768 + 1218) => x"00", (32768 + 1219) => x"00", (32768 + 1220) => x"bc", (32768 + 1221) => x"22", (32768 + 1222) => x"3c", (32768 + 1223) => x"28", (32768 + 1224) => x"a4", (32768 + 1225) => x"89", (32768 + 1226) => x"8a", (32768 + 1227) => x"ab", (32768 + 1228) => x"52", (32768 + 1229) => x"97", (32768 + 1230) => x"51", (32768 + 1231) => x"d1", (32768 + 1232) => x"51", (32768 + 1233) => x"c0", (32768 + 1234) => x"00", (32768 + 1235) => x"00", (32768 + 1236) => x"15", (32768 + 1237) => x"6a", (32768 + 1238) => x"8a", (32768 + 1239) => x"8e", (32768 + 1240) => x"8a", (32768 + 1241) => x"6a", (32768 + 1242) => x"00", (32768 + 1243) => x"64", (32768 + 1244) => x"8a", (32768 + 1245) => x"8e", (32768 + 1246) => x"8a", (32768 + 1247) => x"6a", (32768 + 1248) => x"44", (32768 + 1249) => x"aa", (32768 + 1250) => x"aa", (32768 + 1251) => x"aa", (32768 + 1252) => x"44", (32768 + 1253) => x"00", (32768 + 1254) => x"cc", (32768 + 1255) => x"aa", (32768 + 1256) => x"ca", (32768 + 1257) => x"aa", (32768 + 1258) => x"ac", (32768 + 1259) => x"6e", (32768 + 1260) => x"88", (32768 + 1261) => x"4c", (32768 + 1262) => x"28", (32768 + 1263) => x"ce", (32768 + 1264) => x"00", (32768 + 1265) => x"04", (32768 + 1266) => x"0c", (32768 + 1267) => x"04", (32768 + 1268) => x"04", (32768 + 1269) => x"0e", (32768 + 1270) => x"0c", (32768 + 1271) => x"12", (32768 + 1272) => x"04", (32768 + 1273) => x"08", (32768 + 1274) => x"1e", (32768 + 1275) => x"63", (32768 + 1276) => x"94", (32768 + 1277) => x"94", (32768 + 1278) => x"94", (32768 + 1279) => x"63", (32768 + 1280) => x"38", (32768 + 1281) => x"a5", (32768 + 1282) => x"b8", (32768 + 1283) => x"a0", (32768 + 1284) => x"21", (32768 + 1285) => x"e1", (32768 + 1286) => x"01", (32768 + 1287) => x"c1", (32768 + 1288) => x"20", (32768 + 1289) => x"c1", (32768 + 1290) => x"89", (32768 + 1291) => x"8a", (32768 + 1292) => x"52", (32768 + 1293) => x"22", (32768 + 1294) => x"21", (32768 + 1295) => x"cf", (32768 + 1296) => x"28", (32768 + 1297) => x"2f", (32768 + 1298) => x"28", (32768 + 1299) => x"c8", (32768 + 1300) => x"02", (32768 + 1301) => x"82", (32768 + 1302) => x"02", (32768 + 1303) => x"00", (32768 + 1304) => x"02", (32768 + 1305) => x"ff", (32768 + 1306) => x"80", (32768 + 1307) => x"8f", (32768 + 1308) => x"90", (32768 + 1309) => x"8e", (32768 + 1310) => x"81", (32768 + 1311) => x"9e", (32768 + 1312) => x"80", (32768 + 1313) => x"91", (32768 + 1314) => x"91", (32768 + 1315) => x"9f", (32768 + 1316) => x"91", (32768 + 1317) => x"91", (32768 + 1318) => x"80", (32768 + 1319) => x"ff", (32768 + 1320) => x"00", (32768 + 1321) => x"3c", (32768 + 1322) => x"40", (32768 + 1323) => x"40", (32768 + 1324) => x"40", (32768 + 1325) => x"3c", (32768 + 1326) => x"00", (32768 + 1327) => x"7c", (32768 + 1328) => x"10", (32768 + 1329) => x"10", (32768 + 1330) => x"10", (32768 + 1331) => x"7c", (32768 + 1332) => x"00", (32768 + 1333) => x"ff", (32768 + 1334) => x"00", (32768 + 1335) => x"00", (32768 + 1336) => x"80", (32768 + 1337) => x"00", (32768 + 1338) => x"80", (32768 + 1339) => x"00", (32768 + 1340) => x"00", (32768 + 1341) => x"00", (32768 + 1342) => x"80", (32768 + 1343) => x"00", (32768 + 1344) => x"80", (32768 + 1345) => x"00", (32768 + 1346) => x"00", (32768 + 1347) => x"ff", (32768 + 1348) => x"01", (32768 + 1349) => x"01", (32768 + 1350) => x"01", (32768 + 1351) => x"01", (32768 + 1352) => x"01", (32768 + 1353) => x"01", (32768 + 1354) => x"01", (32768 + 1355) => x"01", (32768 + 1356) => x"01", (32768 + 1357) => x"01", (32768 + 1358) => x"01", (32768 + 1359) => x"01", (32768 + 1360) => x"01", (32768 + 1361) => x"ff", 
                                
                                -- Kaleid by Joseph Weisbecker (RCA)
                                (36864 + 128) => x"00", (36864 + 129) => x"B0", 
                                (36864 + 130) => x"CD", (36864 + 131) => x"E0",
                                (36864 + 132) => x"F0", (36864 + 133) => x"00",
                                (36864 + 134) => x"BE", (36864 + 135) => x"00",
                                (36864 + 136) => x"00", (36864 + 137) => x"20", -- delay
                                (36864 + 138) => x"00",
                                (36864 + 512) => x"60", (36864 + 513) => x"00", (36864 + 514) => x"63", (36864 + 515) => x"80", (36864 + 516) => x"61", (36864 + 517) => x"1f", (36864 + 518) => x"62", (36864 + 519) => x"0f", (36864 + 520) => x"22", (36864 + 521) => x"32", (36864 + 522) => x"a2", (36864 + 523) => x"00", (36864 + 524) => x"f3", (36864 + 525) => x"1e", (36864 + 526) => x"f0", (36864 + 527) => x"0a", (36864 + 528) => x"f0", (36864 + 529) => x"55", (36864 + 530) => x"40", (36864 + 531) => x"00", (36864 + 532) => x"12", (36864 + 533) => x"1c", (36864 + 534) => x"73", (36864 + 535) => x"01", (36864 + 536) => x"33", (36864 + 537) => x"00", (36864 + 538) => x"12", (36864 + 539) => x"08", (36864 + 540) => x"63", (36864 + 541) => x"80", (36864 + 542) => x"a2", (36864 + 543) => x"00", (36864 + 544) => x"f3", (36864 + 545) => x"1e", (36864 + 546) => x"f0", (36864 + 547) => x"65", (36864 + 548) => x"40", (36864 + 549) => x"00", (36864 + 550) => x"12", (36864 + 551) => x"1c", (36864 + 552) => x"73", (36864 + 553) => x"01", (36864 + 554) => x"43", (36864 + 555) => x"00", (36864 + 556) => x"12", (36864 + 557) => x"1c", (36864 + 558) => x"22", (36864 + 559) => x"32", (36864 + 560) => x"12", (36864 + 561) => x"1e", (36864 + 562) => x"40", (36864 + 563) => x"02", (36864 + 564) => x"72", (36864 + 565) => x"ff", (36864 + 566) => x"40", (36864 + 567) => x"04", (36864 + 568) => x"71", (36864 + 569) => x"ff", (36864 + 570) => x"40", (36864 + 571) => x"06", (36864 + 572) => x"71", (36864 + 573) => x"01", (36864 + 574) => x"40", (36864 + 575) => x"08", (36864 + 576) => x"72", (36864 + 577) => x"01", (36864 + 578) => x"a2", (36864 + 579) => x"77", (36864 + 580) => x"6a", (36864 + 581) => x"e0", (36864 + 582) => x"8a", (36864 + 583) => x"12", (36864 + 584) => x"6b", (36864 + 585) => x"1f", (36864 + 586) => x"81", (36864 + 587) => x"b2", (36864 + 588) => x"3a", (36864 + 589) => x"00", (36864 + 590) => x"72", (36864 + 591) => x"01", (36864 + 592) => x"6a", (36864 + 593) => x"f0", (36864 + 594) => x"8a", (36864 + 595) => x"22", (36864 + 596) => x"6b", (36864 + 597) => x"0f", (36864 + 598) => x"82", (36864 + 599) => x"b2", (36864 + 600) => x"3a", (36864 + 601) => x"00", (36864 + 602) => x"71", (36864 + 603) => x"01", (36864 + 604) => x"6b", (36864 + 605) => x"1f", (36864 + 606) => x"81", (36864 + 607) => x"b2", (36864 + 608) => x"d1", (36864 + 609) => x"21", (36864 + 610) => x"8a", (36864 + 611) => x"10", (36864 + 612) => x"6b", (36864 + 613) => x"1f", (36864 + 614) => x"8b", (36864 + 615) => x"25", (36864 + 616) => x"da", (36864 + 617) => x"b1", (36864 + 618) => x"6a", (36864 + 619) => x"3f", (36864 + 620) => x"8a", (36864 + 621) => x"15", (36864 + 622) => x"da", (36864 + 623) => x"b1", (36864 + 624) => x"8b", (36864 + 625) => x"20", (36864 + 626) => x"da", (36864 + 627) => x"b1", (36864 + 628) => x"00", (36864 + 629) => x"ee", (36864 + 630) => x"01", (36864 + 631) => x"80", 
                                
                                -- Merlin by David Winter
                                (40960 + 128) => x"00", (40960 + 129) => x"00", 
                                (40960 + 130) => x"CB", (40960 + 131) => x"0F",
                                (40960 + 132) => x"E0", (40960 + 133) => x"00",
                                (40960 + 134) => x"BE", (40960 + 135) => x"00",
                                (40960 + 136) => x"00", (40960 + 137) => x"30", -- delay
                                (40960 + 138) => x"00",
                                (40960 + 512) => x"12", (40960 + 513) => x"19", (40960 + 514) => x"20", (40960 + 515) => x"4d", (40960 + 516) => x"45", (40960 + 517) => x"52", (40960 + 518) => x"4c", (40960 + 519) => x"49", (40960 + 520) => x"4e", (40960 + 521) => x"20", (40960 + 522) => x"42", (40960 + 523) => x"79", (40960 + 524) => x"20", (40960 + 525) => x"44", (40960 + 526) => x"61", (40960 + 527) => x"76", (40960 + 528) => x"69", (40960 + 529) => x"64", (40960 + 530) => x"20", (40960 + 531) => x"57", (40960 + 532) => x"49", (40960 + 533) => x"4e", (40960 + 534) => x"54", (40960 + 535) => x"45", (40960 + 536) => x"52", (40960 + 537) => x"22", (40960 + 538) => x"f9", (40960 + 539) => x"a3", (40960 + 540) => x"1d", (40960 + 541) => x"60", (40960 + 542) => x"10", (40960 + 543) => x"61", (40960 + 544) => x"00", (40960 + 545) => x"22", (40960 + 546) => x"cb", (40960 + 547) => x"a3", (40960 + 548) => x"31", (40960 + 549) => x"60", (40960 + 550) => x"0b", (40960 + 551) => x"61", (40960 + 552) => x"1b", (40960 + 553) => x"22", (40960 + 554) => x"cb", (40960 + 555) => x"64", (40960 + 556) => x"04", (40960 + 557) => x"22", (40960 + 558) => x"df", (40960 + 559) => x"65", (40960 + 560) => x"00", (40960 + 561) => x"62", (40960 + 562) => x"28", (40960 + 563) => x"22", (40960 + 564) => x"c1", (40960 + 565) => x"c2", (40960 + 566) => x"03", (40960 + 567) => x"80", (40960 + 568) => x"20", (40960 + 569) => x"a3", (40960 + 570) => x"59", (40960 + 571) => x"f5", (40960 + 572) => x"1e", (40960 + 573) => x"f0", (40960 + 574) => x"55", (40960 + 575) => x"60", (40960 + 576) => x"17", (40960 + 577) => x"61", (40960 + 578) => x"08", (40960 + 579) => x"63", (40960 + 580) => x"01", (40960 + 581) => x"83", (40960 + 582) => x"22", (40960 + 583) => x"33", (40960 + 584) => x"00", (40960 + 585) => x"70", (40960 + 586) => x"0a", (40960 + 587) => x"63", (40960 + 588) => x"02", (40960 + 589) => x"83", (40960 + 590) => x"22", (40960 + 591) => x"33", (40960 + 592) => x"00", (40960 + 593) => x"71", (40960 + 594) => x"0a", (40960 + 595) => x"a3", (40960 + 596) => x"17", (40960 + 597) => x"d0", (40960 + 598) => x"16", (40960 + 599) => x"62", (40960 + 600) => x"14", (40960 + 601) => x"22", (40960 + 602) => x"c1", (40960 + 603) => x"d0", (40960 + 604) => x"16", (40960 + 605) => x"62", (40960 + 606) => x"05", (40960 + 607) => x"22", (40960 + 608) => x"c1", (40960 + 609) => x"75", (40960 + 610) => x"01", (40960 + 611) => x"54", (40960 + 612) => x"50", (40960 + 613) => x"12", (40960 + 614) => x"35", (40960 + 615) => x"65", (40960 + 616) => x"00", (40960 + 617) => x"60", (40960 + 618) => x"17", (40960 + 619) => x"61", (40960 + 620) => x"08", (40960 + 621) => x"a3", (40960 + 622) => x"17", (40960 + 623) => x"f3", (40960 + 624) => x"0a", (40960 + 625) => x"33", (40960 + 626) => x"04", (40960 + 627) => x"12", (40960 + 628) => x"79", (40960 + 629) => x"63", (40960 + 630) => x"00", (40960 + 631) => x"12", (40960 + 632) => x"97", (40960 + 633) => x"33", (40960 + 634) => x"05", (40960 + 635) => x"12", (40960 + 636) => x"83", (40960 + 637) => x"70", (40960 + 638) => x"0a", (40960 + 639) => x"63", (40960 + 640) => x"01", (40960 + 641) => x"12", (40960 + 642) => x"97", (40960 + 643) => x"33", (40960 + 644) => x"07", (40960 + 645) => x"12", (40960 + 646) => x"8d", (40960 + 647) => x"71", (40960 + 648) => x"0a", (40960 + 649) => x"63", (40960 + 650) => x"02", (40960 + 651) => x"12", (40960 + 652) => x"97", (40960 + 653) => x"33", (40960 + 654) => x"08", (40960 + 655) => x"12", (40960 + 656) => x"69", (40960 + 657) => x"70", (40960 + 658) => x"0a", (40960 + 659) => x"71", (40960 + 660) => x"0a", (40960 + 661) => x"63", (40960 + 662) => x"03", (40960 + 663) => x"d0", (40960 + 664) => x"16", (40960 + 665) => x"62", (40960 + 666) => x"14", (40960 + 667) => x"22", (40960 + 668) => x"c1", (40960 + 669) => x"d0", (40960 + 670) => x"16", (40960 + 671) => x"a3", (40960 + 672) => x"59", (40960 + 673) => x"f5", (40960 + 674) => x"1e", (40960 + 675) => x"f0", (40960 + 676) => x"65", (40960 + 677) => x"75", (40960 + 678) => x"01", (40960 + 679) => x"50", (40960 + 680) => x"30", (40960 + 681) => x"12", (40960 + 682) => x"b5", (40960 + 683) => x"55", (40960 + 684) => x"40", (40960 + 685) => x"12", (40960 + 686) => x"69", (40960 + 687) => x"22", (40960 + 688) => x"df", (40960 + 689) => x"74", (40960 + 690) => x"01", (40960 + 691) => x"12", (40960 + 692) => x"2d", (40960 + 693) => x"22", (40960 + 694) => x"f9", (40960 + 695) => x"a3", (40960 + 696) => x"45", (40960 + 697) => x"60", (40960 + 698) => x"10", (40960 + 699) => x"61", (40960 + 700) => x"0e", (40960 + 701) => x"22", (40960 + 702) => x"cb", (40960 + 703) => x"12", (40960 + 704) => x"bf", (40960 + 705) => x"f2", (40960 + 706) => x"15", (40960 + 707) => x"f2", (40960 + 708) => x"07", (40960 + 709) => x"32", (40960 + 710) => x"00", (40960 + 711) => x"12", (40960 + 712) => x"c3", (40960 + 713) => x"00", (40960 + 714) => x"ee", (40960 + 715) => x"83", (40960 + 716) => x"00", (40960 + 717) => x"62", (40960 + 718) => x"05", (40960 + 719) => x"d0", (40960 + 720) => x"15", (40960 + 721) => x"f2", (40960 + 722) => x"1e", (40960 + 723) => x"70", (40960 + 724) => x"08", (40960 + 725) => x"85", (40960 + 726) => x"30", (40960 + 727) => x"75", (40960 + 728) => x"20", (40960 + 729) => x"50", (40960 + 730) => x"50", (40960 + 731) => x"12", (40960 + 732) => x"cf", (40960 + 733) => x"00", (40960 + 734) => x"ee", (40960 + 735) => x"a3", (40960 + 736) => x"59", (40960 + 737) => x"83", (40960 + 738) => x"40", (40960 + 739) => x"73", (40960 + 740) => x"fd", (40960 + 741) => x"f3", (40960 + 742) => x"33", (40960 + 743) => x"f2", (40960 + 744) => x"65", (40960 + 745) => x"f1", (40960 + 746) => x"29", (40960 + 747) => x"60", (40960 + 748) => x"2b", (40960 + 749) => x"63", (40960 + 750) => x"1b", (40960 + 751) => x"d0", (40960 + 752) => x"35", (40960 + 753) => x"70", (40960 + 754) => x"05", (40960 + 755) => x"f2", (40960 + 756) => x"29", (40960 + 757) => x"d0", (40960 + 758) => x"35", (40960 + 759) => x"00", (40960 + 760) => x"ee", (40960 + 761) => x"a3", (40960 + 762) => x"0f", (40960 + 763) => x"60", (40960 + 764) => x"17", (40960 + 765) => x"61", (40960 + 766) => x"07", (40960 + 767) => x"d0", (40960 + 768) => x"18", (40960 + 769) => x"70", (40960 + 770) => x"0a", (40960 + 771) => x"d0", (40960 + 772) => x"18", (40960 + 773) => x"71", (40960 + 774) => x"0a", (40960 + 775) => x"d0", (40960 + 776) => x"18", (40960 + 777) => x"70", (40960 + 778) => x"f6", (40960 + 779) => x"d0", (40960 + 780) => x"18", (40960 + 781) => x"00", (40960 + 782) => x"ee", (40960 + 783) => x"ff", (40960 + 784) => x"81", (40960 + 785) => x"81", (40960 + 786) => x"81", (40960 + 787) => x"81", (40960 + 788) => x"81", (40960 + 789) => x"81", (40960 + 790) => x"ff", (40960 + 791) => x"7e", (40960 + 792) => x"7e", (40960 + 793) => x"7e", (40960 + 794) => x"7e", (40960 + 795) => x"7e", (40960 + 796) => x"7e", (40960 + 797) => x"db", (40960 + 798) => x"aa", (40960 + 799) => x"8b", (40960 + 800) => x"cb", (40960 + 801) => x"cb", (40960 + 802) => x"ef", (40960 + 803) => x"08", (40960 + 804) => x"8f", (40960 + 805) => x"0d", (40960 + 806) => x"ec", (40960 + 807) => x"a0", (40960 + 808) => x"a0", (40960 + 809) => x"b0", (40960 + 810) => x"30", (40960 + 811) => x"be", (40960 + 812) => x"5f", (40960 + 813) => x"51", (40960 + 814) => x"51", (40960 + 815) => x"d9", (40960 + 816) => x"d9", (40960 + 817) => x"83", (40960 + 818) => x"82", (40960 + 819) => x"83", (40960 + 820) => x"82", (40960 + 821) => x"fb", (40960 + 822) => x"e8", (40960 + 823) => x"08", (40960 + 824) => x"88", (40960 + 825) => x"05", (40960 + 826) => x"e2", (40960 + 827) => x"be", (40960 + 828) => x"a0", (40960 + 829) => x"b8", (40960 + 830) => x"20", (40960 + 831) => x"3e", (40960 + 832) => x"80", (40960 + 833) => x"80", (40960 + 834) => x"80", (40960 + 835) => x"80", (40960 + 836) => x"f8", (40960 + 837) => x"f7", (40960 + 838) => x"85", (40960 + 839) => x"b7", (40960 + 840) => x"95", (40960 + 841) => x"f5", (40960 + 842) => x"76", (40960 + 843) => x"54", (40960 + 844) => x"56", (40960 + 845) => x"54", (40960 + 846) => x"56", (40960 + 847) => x"3a", (40960 + 848) => x"2a", (40960 + 849) => x"2a", (40960 + 850) => x"2a", (40960 + 851) => x"39", (40960 + 852) => x"b6", (40960 + 853) => x"a5", (40960 + 854) => x"b6", (40960 + 855) => x"a5", (40960 + 856) => x"35", (40960 + 857) => x"00", 
                                
                                -- Missile by David Winter 
                                (45056 + 128) => x"0F", (45056 + 129) => x"00", 
                                (45056 + 130) => x"C0", (45056 + 131) => x"00",
                                (45056 + 132) => x"D0", (45056 + 133) => x"00",
                                (45056 + 134) => x"BE", (45056 + 135) => x"00",
                                (45056 + 136) => x"00", (45056 + 137) => x"30", -- delay
                                (45056 + 138) => x"00",
                                (45056 + 512) => x"12", (45056 + 513) => x"19", (45056 + 514) => x"4d", (45056 + 515) => x"49", (45056 + 516) => x"53", (45056 + 517) => x"53", (45056 + 518) => x"49", (45056 + 519) => x"4c", (45056 + 520) => x"45", (45056 + 521) => x"20", (45056 + 522) => x"62", (45056 + 523) => x"79", (45056 + 524) => x"20", (45056 + 525) => x"44", (45056 + 526) => x"61", (45056 + 527) => x"76", (45056 + 528) => x"69", (45056 + 529) => x"64", (45056 + 530) => x"20", (45056 + 531) => x"57", (45056 + 532) => x"49", (45056 + 533) => x"4e", (45056 + 534) => x"54", (45056 + 535) => x"45", (45056 + 536) => x"52", (45056 + 537) => x"6c", (45056 + 538) => x"0c", (45056 + 539) => x"60", (45056 + 540) => x"00", (45056 + 541) => x"61", (45056 + 542) => x"00", (45056 + 543) => x"65", (45056 + 544) => x"08", (45056 + 545) => x"66", (45056 + 546) => x"0a", (45056 + 547) => x"67", (45056 + 548) => x"00", (45056 + 549) => x"6e", (45056 + 550) => x"01", (45056 + 551) => x"a2", (45056 + 552) => x"ad", (45056 + 553) => x"d0", (45056 + 554) => x"14", (45056 + 555) => x"70", (45056 + 556) => x"08", (45056 + 557) => x"30", (45056 + 558) => x"40", (45056 + 559) => x"12", (45056 + 560) => x"29", (45056 + 561) => x"60", (45056 + 562) => x"00", (45056 + 563) => x"61", (45056 + 564) => x"1c", (45056 + 565) => x"a2", (45056 + 566) => x"b0", (45056 + 567) => x"d0", (45056 + 568) => x"14", (45056 + 569) => x"a2", (45056 + 570) => x"b0", (45056 + 571) => x"d0", (45056 + 572) => x"14", (45056 + 573) => x"3e", (45056 + 574) => x"01", (45056 + 575) => x"12", (45056 + 576) => x"49", (45056 + 577) => x"70", (45056 + 578) => x"04", (45056 + 579) => x"40", (45056 + 580) => x"38", (45056 + 581) => x"6e", (45056 + 582) => x"00", (45056 + 583) => x"12", (45056 + 584) => x"4f", (45056 + 585) => x"70", (45056 + 586) => x"fc", (45056 + 587) => x"40", (45056 + 588) => x"00", (45056 + 589) => x"6e", (45056 + 590) => x"01", (45056 + 591) => x"d0", (45056 + 592) => x"14", (45056 + 593) => x"fc", (45056 + 594) => x"15", (45056 + 595) => x"fb", (45056 + 596) => x"07", (45056 + 597) => x"3b", (45056 + 598) => x"00", (45056 + 599) => x"12", (45056 + 600) => x"53", (45056 + 601) => x"62", (45056 + 602) => x"08", (45056 + 603) => x"e2", (45056 + 604) => x"9e", (45056 + 605) => x"12", (45056 + 606) => x"95", (45056 + 607) => x"3c", (45056 + 608) => x"00", (45056 + 609) => x"7c", (45056 + 610) => x"fe", (45056 + 611) => x"63", (45056 + 612) => x"1b", (45056 + 613) => x"82", (45056 + 614) => x"00", (45056 + 615) => x"a2", (45056 + 616) => x"b0", (45056 + 617) => x"d2", (45056 + 618) => x"31", (45056 + 619) => x"64", (45056 + 620) => x"00", (45056 + 621) => x"d2", (45056 + 622) => x"31", (45056 + 623) => x"73", (45056 + 624) => x"ff", (45056 + 625) => x"d2", (45056 + 626) => x"31", (45056 + 627) => x"3f", (45056 + 628) => x"00", (45056 + 629) => x"64", (45056 + 630) => x"01", (45056 + 631) => x"33", (45056 + 632) => x"03", (45056 + 633) => x"12", (45056 + 634) => x"6d", (45056 + 635) => x"d2", (45056 + 636) => x"31", (45056 + 637) => x"34", (45056 + 638) => x"01", (45056 + 639) => x"12", (45056 + 640) => x"91", (45056 + 641) => x"77", (45056 + 642) => x"05", (45056 + 643) => x"75", (45056 + 644) => x"ff", (45056 + 645) => x"82", (45056 + 646) => x"00", (45056 + 647) => x"63", (45056 + 648) => x"00", (45056 + 649) => x"a2", (45056 + 650) => x"ad", (45056 + 651) => x"d2", (45056 + 652) => x"34", (45056 + 653) => x"45", (45056 + 654) => x"00", (45056 + 655) => x"12", (45056 + 656) => x"97", (45056 + 657) => x"76", (45056 + 658) => x"ff", (45056 + 659) => x"36", (45056 + 660) => x"00", (45056 + 661) => x"12", (45056 + 662) => x"39", (45056 + 663) => x"a2", (45056 + 664) => x"b4", (45056 + 665) => x"f7", (45056 + 666) => x"33", (45056 + 667) => x"f2", (45056 + 668) => x"65", (45056 + 669) => x"63", (45056 + 670) => x"1b", (45056 + 671) => x"64", (45056 + 672) => x"0d", (45056 + 673) => x"f1", (45056 + 674) => x"29", (45056 + 675) => x"d3", (45056 + 676) => x"45", (45056 + 677) => x"73", (45056 + 678) => x"05", (45056 + 679) => x"f2", (45056 + 680) => x"29", (45056 + 681) => x"d3", (45056 + 682) => x"45", (45056 + 683) => x"12", (45056 + 684) => x"ab", (45056 + 685) => x"10", (45056 + 686) => x"38", (45056 + 687) => x"38", (45056 + 688) => x"10", (45056 + 689) => x"38", (45056 + 690) => x"7c", (45056 + 691) => x"fe", 
                                
                                -- Puzzle by Joseph Weisbecker (RCA)
                                (49152 + 128) => x"00", (49152 + 129) => x"B0", 
                                (49152 + 130) => x"C0", (49152 + 131) => x"E0",
                                (49152 + 132) => x"F0", (49152 + 133) => x"00",
                                (49152 + 134) => x"BE", (49152 + 135) => x"00",
                                (49152 + 136) => x"00", (49152 + 137) => x"30", -- delay
                                (49152 + 138) => x"00",
                                (49152 + 512) => x"6a", (49152 + 513) => x"12", (49152 + 514) => x"6b", (49152 + 515) => x"01", (49152 + 516) => x"61", (49152 + 517) => x"10", (49152 + 518) => x"62", (49152 + 519) => x"00", (49152 + 520) => x"60", (49152 + 521) => x"00", (49152 + 522) => x"a2", (49152 + 523) => x"b0", (49152 + 524) => x"d1", (49152 + 525) => x"27", (49152 + 526) => x"f0", (49152 + 527) => x"29", (49152 + 528) => x"30", (49152 + 529) => x"00", (49152 + 530) => x"da", (49152 + 531) => x"b5", (49152 + 532) => x"71", (49152 + 533) => x"08", (49152 + 534) => x"7a", (49152 + 535) => x"08", (49152 + 536) => x"31", (49152 + 537) => x"30", (49152 + 538) => x"12", (49152 + 539) => x"24", (49152 + 540) => x"61", (49152 + 541) => x"10", (49152 + 542) => x"72", (49152 + 543) => x"08", (49152 + 544) => x"6a", (49152 + 545) => x"12", (49152 + 546) => x"7b", (49152 + 547) => x"08", (49152 + 548) => x"a3", (49152 + 549) => x"00", (49152 + 550) => x"f0", (49152 + 551) => x"1e", (49152 + 552) => x"f0", (49152 + 553) => x"55", (49152 + 554) => x"70", (49152 + 555) => x"01", (49152 + 556) => x"30", (49152 + 557) => x"10", (49152 + 558) => x"12", (49152 + 559) => x"0a", (49152 + 560) => x"6a", (49152 + 561) => x"12", (49152 + 562) => x"6b", (49152 + 563) => x"01", (49152 + 564) => x"6c", (49152 + 565) => x"00", (49152 + 566) => x"62", (49152 + 567) => x"ff", (49152 + 568) => x"c0", (49152 + 569) => x"06", (49152 + 570) => x"70", (49152 + 571) => x"02", (49152 + 572) => x"22", (49152 + 573) => x"52", (49152 + 574) => x"72", (49152 + 575) => x"ff", (49152 + 576) => x"32", (49152 + 577) => x"00", (49152 + 578) => x"12", (49152 + 579) => x"38", (49152 + 580) => x"6e", (49152 + 581) => x"00", (49152 + 582) => x"6e", (49152 + 583) => x"00", (49152 + 584) => x"f0", (49152 + 585) => x"0a", (49152 + 586) => x"22", (49152 + 587) => x"52", (49152 + 588) => x"7e", (49152 + 589) => x"01", (49152 + 590) => x"7e", (49152 + 591) => x"01", (49152 + 592) => x"12", (49152 + 593) => x"48", (49152 + 594) => x"84", (49152 + 595) => x"a0", (49152 + 596) => x"85", (49152 + 597) => x"b0", (49152 + 598) => x"86", (49152 + 599) => x"c0", (49152 + 600) => x"30", (49152 + 601) => x"02", (49152 + 602) => x"12", (49152 + 603) => x"64", (49152 + 604) => x"45", (49152 + 605) => x"01", (49152 + 606) => x"12", (49152 + 607) => x"64", (49152 + 608) => x"75", (49152 + 609) => x"f8", (49152 + 610) => x"76", (49152 + 611) => x"fc", (49152 + 612) => x"30", (49152 + 613) => x"08", (49152 + 614) => x"12", (49152 + 615) => x"70", (49152 + 616) => x"45", (49152 + 617) => x"19", (49152 + 618) => x"12", (49152 + 619) => x"70", (49152 + 620) => x"75", (49152 + 621) => x"08", (49152 + 622) => x"76", (49152 + 623) => x"04", (49152 + 624) => x"30", (49152 + 625) => x"06", (49152 + 626) => x"12", (49152 + 627) => x"7c", (49152 + 628) => x"44", (49152 + 629) => x"12", (49152 + 630) => x"12", (49152 + 631) => x"7c", (49152 + 632) => x"74", (49152 + 633) => x"f8", (49152 + 634) => x"76", (49152 + 635) => x"ff", (49152 + 636) => x"30", (49152 + 637) => x"04", (49152 + 638) => x"12", (49152 + 639) => x"88", (49152 + 640) => x"44", (49152 + 641) => x"2a", (49152 + 642) => x"12", (49152 + 643) => x"88", (49152 + 644) => x"74", (49152 + 645) => x"08", (49152 + 646) => x"76", (49152 + 647) => x"01", (49152 + 648) => x"a3", (49152 + 649) => x"00", (49152 + 650) => x"f6", (49152 + 651) => x"1e", (49152 + 652) => x"f0", (49152 + 653) => x"65", (49152 + 654) => x"81", (49152 + 655) => x"00", (49152 + 656) => x"60", (49152 + 657) => x"00", (49152 + 658) => x"a3", (49152 + 659) => x"00", (49152 + 660) => x"f6", (49152 + 661) => x"1e", (49152 + 662) => x"f0", (49152 + 663) => x"55", (49152 + 664) => x"a3", (49152 + 665) => x"00", (49152 + 666) => x"fc", (49152 + 667) => x"1e", (49152 + 668) => x"80", (49152 + 669) => x"10", (49152 + 670) => x"f0", (49152 + 671) => x"55", (49152 + 672) => x"f1", (49152 + 673) => x"29", (49152 + 674) => x"d4", (49152 + 675) => x"55", (49152 + 676) => x"da", (49152 + 677) => x"b5", (49152 + 678) => x"8a", (49152 + 679) => x"40", (49152 + 680) => x"8b", (49152 + 681) => x"50", (49152 + 682) => x"8c", (49152 + 683) => x"60", (49152 + 684) => x"00", (49152 + 685) => x"ee", (49152 + 686) => x"ee", (49152 + 687) => x"5e", (49152 + 688) => x"fe", (49152 + 689) => x"fe", (49152 + 690) => x"fe", (49152 + 691) => x"fe", (49152 + 692) => x"fe", (49152 + 693) => x"fe", (49152 + 694) => x"fe", (49152 + 695) => x"fe", 
                                
                                -- Tank by Joseph Weisbecker (RCA)
                                (53248 + 128) => x"00", (53248 + 129) => x"B0", 
                                (53248 + 130) => x"CD", (53248 + 131) => x"E0",
                                (53248 + 132) => x"F0", (53248 + 133) => x"00",
                                (53248 + 134) => x"BE", (53248 + 135) => x"00",
                                (53248 + 136) => x"00", (53248 + 137) => x"30", -- delay
                                (53248 + 138) => x"00",
                                (53248 + 512) => x"12", (53248 + 513) => x"30", (53248 + 514) => x"76", (53248 + 515) => x"fb", (53248 + 516) => x"60", (53248 + 517) => x"20", (53248 + 518) => x"80", (53248 + 519) => x"65", (53248 + 520) => x"4f", (53248 + 521) => x"00", (53248 + 522) => x"66", (53248 + 523) => x"00", (53248 + 524) => x"13", (53248 + 525) => x"84", (53248 + 526) => x"00", (53248 + 527) => x"ff", (53248 + 528) => x"00", (53248 + 529) => x"00", (53248 + 530) => x"00", (53248 + 531) => x"01", (53248 + 532) => x"00", (53248 + 533) => x"0c", (53248 + 534) => x"0a", (53248 + 535) => x"00", (53248 + 536) => x"19", (53248 + 537) => x"02", (53248 + 538) => x"04", (53248 + 539) => x"06", (53248 + 540) => x"08", (53248 + 541) => x"02", (53248 + 542) => x"02", (53248 + 543) => x"03", (53248 + 544) => x"2c", (53248 + 545) => x"00", (53248 + 546) => x"0f", (53248 + 547) => x"00", (53248 + 548) => x"02", (53248 + 549) => x"05", (53248 + 550) => x"2e", (53248 + 551) => x"08", (53248 + 552) => x"00", (53248 + 553) => x"00", (53248 + 554) => x"02", (53248 + 555) => x"05", (53248 + 556) => x"00", (53248 + 557) => x"00", (53248 + 558) => x"00", (53248 + 559) => x"00", (53248 + 560) => x"6e", (53248 + 561) => x"00", (53248 + 562) => x"6d", (53248 + 563) => x"a0", (53248 + 564) => x"6a", (53248 + 565) => x"08", (53248 + 566) => x"69", (53248 + 567) => x"06", (53248 + 568) => x"68", (53248 + 569) => x"04", (53248 + 570) => x"67", (53248 + 571) => x"02", (53248 + 572) => x"66", (53248 + 573) => x"19", (53248 + 574) => x"64", (53248 + 575) => x"10", (53248 + 576) => x"63", (53248 + 577) => x"0c", (53248 + 578) => x"62", (53248 + 579) => x"00", (53248 + 580) => x"61", (53248 + 581) => x"06", (53248 + 582) => x"a2", (53248 + 583) => x"12", (53248 + 584) => x"fa", (53248 + 585) => x"55", (53248 + 586) => x"23", (53248 + 587) => x"d4", (53248 + 588) => x"60", (53248 + 589) => x"40", (53248 + 590) => x"f0", (53248 + 591) => x"15", (53248 + 592) => x"f0", (53248 + 593) => x"07", (53248 + 594) => x"30", (53248 + 595) => x"00", (53248 + 596) => x"12", (53248 + 597) => x"50", (53248 + 598) => x"23", (53248 + 599) => x"d4", (53248 + 600) => x"23", (53248 + 601) => x"0a", (53248 + 602) => x"23", (53248 + 603) => x"62", (53248 + 604) => x"a2", (53248 + 605) => x"12", (53248 + 606) => x"f5", (53248 + 607) => x"65", (53248 + 608) => x"22", (53248 + 609) => x"ae", (53248 + 610) => x"22", (53248 + 611) => x"c6", (53248 + 612) => x"22", (53248 + 613) => x"ec", (53248 + 614) => x"3f", (53248 + 615) => x"01", (53248 + 616) => x"23", (53248 + 617) => x"14", (53248 + 618) => x"3f", (53248 + 619) => x"01", (53248 + 620) => x"22", (53248 + 621) => x"ec", (53248 + 622) => x"3f", (53248 + 623) => x"01", (53248 + 624) => x"22", (53248 + 625) => x"ec", (53248 + 626) => x"3f", (53248 + 627) => x"01", (53248 + 628) => x"22", (53248 + 629) => x"7c", (53248 + 630) => x"4f", (53248 + 631) => x"01", (53248 + 632) => x"13", (53248 + 633) => x"66", (53248 + 634) => x"12", (53248 + 635) => x"62", (53248 + 636) => x"a2", (53248 + 637) => x"12", (53248 + 638) => x"f5", (53248 + 639) => x"65", (53248 + 640) => x"46", (53248 + 641) => x"00", (53248 + 642) => x"35", (53248 + 643) => x"00", (53248 + 644) => x"12", (53248 + 645) => x"88", (53248 + 646) => x"13", (53248 + 647) => x"8c", (53248 + 648) => x"e7", (53248 + 649) => x"a1", (53248 + 650) => x"62", (53248 + 651) => x"09", (53248 + 652) => x"e8", (53248 + 653) => x"a1", (53248 + 654) => x"62", (53248 + 655) => x"04", (53248 + 656) => x"e9", (53248 + 657) => x"a1", (53248 + 658) => x"62", (53248 + 659) => x"06", (53248 + 660) => x"ea", (53248 + 661) => x"a1", (53248 + 662) => x"62", (53248 + 663) => x"01", (53248 + 664) => x"42", (53248 + 665) => x"00", (53248 + 666) => x"00", (53248 + 667) => x"ee", (53248 + 668) => x"22", (53248 + 669) => x"ae", (53248 + 670) => x"81", (53248 + 671) => x"20", (53248 + 672) => x"23", (53248 + 673) => x"9a", (53248 + 674) => x"23", (53248 + 675) => x"ac", (53248 + 676) => x"6c", (53248 + 677) => x"01", (53248 + 678) => x"62", (53248 + 679) => x"00", (53248 + 680) => x"6f", (53248 + 681) => x"00", (53248 + 682) => x"a2", (53248 + 683) => x"12", (53248 + 684) => x"f5", (53248 + 685) => x"55", (53248 + 686) => x"a3", (53248 + 687) => x"ff", (53248 + 688) => x"41", (53248 + 689) => x"01", (53248 + 690) => x"60", (53248 + 691) => x"00", (53248 + 692) => x"41", (53248 + 693) => x"04", (53248 + 694) => x"60", (53248 + 695) => x"13", (53248 + 696) => x"41", (53248 + 697) => x"06", (53248 + 698) => x"60", (53248 + 699) => x"0d", (53248 + 700) => x"41", (53248 + 701) => x"09", (53248 + 702) => x"60", (53248 + 703) => x"06", (53248 + 704) => x"f0", (53248 + 705) => x"1e", (53248 + 706) => x"d3", (53248 + 707) => x"47", (53248 + 708) => x"00", (53248 + 709) => x"ee", (53248 + 710) => x"60", (53248 + 711) => x"05", (53248 + 712) => x"e0", (53248 + 713) => x"9e", (53248 + 714) => x"00", (53248 + 715) => x"ee", (53248 + 716) => x"45", (53248 + 717) => x"0f", (53248 + 718) => x"00", (53248 + 719) => x"ee", (53248 + 720) => x"65", (53248 + 721) => x"0f", (53248 + 722) => x"76", (53248 + 723) => x"ff", (53248 + 724) => x"a2", (53248 + 725) => x"12", (53248 + 726) => x"f5", (53248 + 727) => x"55", (53248 + 728) => x"74", (53248 + 729) => x"03", (53248 + 730) => x"73", (53248 + 731) => x"03", (53248 + 732) => x"23", (53248 + 733) => x"9a", (53248 + 734) => x"23", (53248 + 735) => x"9a", (53248 + 736) => x"23", (53248 + 737) => x"9a", (53248 + 738) => x"a2", (53248 + 739) => x"23", (53248 + 740) => x"f5", (53248 + 741) => x"55", (53248 + 742) => x"a4", (53248 + 743) => x"19", (53248 + 744) => x"d3", (53248 + 745) => x"41", (53248 + 746) => x"00", (53248 + 747) => x"ee", (53248 + 748) => x"a2", (53248 + 749) => x"23", (53248 + 750) => x"f5", (53248 + 751) => x"65", (53248 + 752) => x"45", (53248 + 753) => x"00", (53248 + 754) => x"00", (53248 + 755) => x"ee", (53248 + 756) => x"a4", (53248 + 757) => x"19", (53248 + 758) => x"d3", (53248 + 759) => x"41", (53248 + 760) => x"23", (53248 + 761) => x"9a", (53248 + 762) => x"6c", (53248 + 763) => x"02", (53248 + 764) => x"23", (53248 + 765) => x"be", (53248 + 766) => x"4b", (53248 + 767) => x"bb", (53248 + 768) => x"13", (53248 + 769) => x"0a", (53248 + 770) => x"d3", (53248 + 771) => x"41", (53248 + 772) => x"a2", (53248 + 773) => x"23", (53248 + 774) => x"f5", (53248 + 775) => x"55", (53248 + 776) => x"00", (53248 + 777) => x"ee", (53248 + 778) => x"65", (53248 + 779) => x"00", (53248 + 780) => x"60", (53248 + 781) => x"00", (53248 + 782) => x"a2", (53248 + 783) => x"17", (53248 + 784) => x"f0", (53248 + 785) => x"55", (53248 + 786) => x"13", (53248 + 787) => x"04", (53248 + 788) => x"a2", (53248 + 789) => x"1d", (53248 + 790) => x"f5", (53248 + 791) => x"65", (53248 + 792) => x"35", (53248 + 793) => x"0f", (53248 + 794) => x"13", (53248 + 795) => x"44", (53248 + 796) => x"a4", (53248 + 797) => x"1a", (53248 + 798) => x"d3", (53248 + 799) => x"45", (53248 + 800) => x"32", (53248 + 801) => x"00", (53248 + 802) => x"13", (53248 + 803) => x"32", (53248 + 804) => x"c1", (53248 + 805) => x"03", (53248 + 806) => x"a2", (53248 + 807) => x"19", (53248 + 808) => x"f1", (53248 + 809) => x"1e", (53248 + 810) => x"f0", (53248 + 811) => x"65", (53248 + 812) => x"81", (53248 + 813) => x"00", (53248 + 814) => x"c2", (53248 + 815) => x"0f", (53248 + 816) => x"72", (53248 + 817) => x"01", (53248 + 818) => x"23", (53248 + 819) => x"9a", (53248 + 820) => x"a4", (53248 + 821) => x"1a", (53248 + 822) => x"6c", (53248 + 823) => x"03", (53248 + 824) => x"72", (53248 + 825) => x"ff", (53248 + 826) => x"6f", (53248 + 827) => x"00", (53248 + 828) => x"d3", (53248 + 829) => x"45", (53248 + 830) => x"a2", (53248 + 831) => x"1d", (53248 + 832) => x"f5", (53248 + 833) => x"55", (53248 + 834) => x"00", (53248 + 835) => x"ee", (53248 + 836) => x"c4", (53248 + 837) => x"07", (53248 + 838) => x"a4", (53248 + 839) => x"1f", (53248 + 840) => x"f4", (53248 + 841) => x"1e", (53248 + 842) => x"f0", (53248 + 843) => x"65", (53248 + 844) => x"83", (53248 + 845) => x"00", (53248 + 846) => x"a4", (53248 + 847) => x"27", (53248 + 848) => x"f4", (53248 + 849) => x"1e", (53248 + 850) => x"f0", (53248 + 851) => x"65", (53248 + 852) => x"84", (53248 + 853) => x"00", (53248 + 854) => x"a4", (53248 + 855) => x"1a", (53248 + 856) => x"d3", (53248 + 857) => x"45", (53248 + 858) => x"60", (53248 + 859) => x"20", (53248 + 860) => x"f0", (53248 + 861) => x"18", (53248 + 862) => x"65", (53248 + 863) => x"0f", (53248 + 864) => x"13", (53248 + 865) => x"3e", (53248 + 866) => x"65", (53248 + 867) => x"00", (53248 + 868) => x"13", (53248 + 869) => x"3e", (53248 + 870) => x"4c", (53248 + 871) => x"01", (53248 + 872) => x"12", (53248 + 873) => x"02", (53248 + 874) => x"4c", (53248 + 875) => x"02", (53248 + 876) => x"13", (53248 + 877) => x"82", (53248 + 878) => x"a2", (53248 + 879) => x"23", (53248 + 880) => x"f5", (53248 + 881) => x"65", (53248 + 882) => x"45", (53248 + 883) => x"00", (53248 + 884) => x"12", (53248 + 885) => x"02", (53248 + 886) => x"a4", (53248 + 887) => x"19", (53248 + 888) => x"d3", (53248 + 889) => x"41", (53248 + 890) => x"6f", (53248 + 891) => x"00", (53248 + 892) => x"d3", (53248 + 893) => x"41", (53248 + 894) => x"3f", (53248 + 895) => x"01", (53248 + 896) => x"12", (53248 + 897) => x"02", (53248 + 898) => x"7e", (53248 + 899) => x"0a", (53248 + 900) => x"60", (53248 + 901) => x"40", (53248 + 902) => x"f0", (53248 + 903) => x"18", (53248 + 904) => x"00", (53248 + 905) => x"e0", (53248 + 906) => x"12", (53248 + 907) => x"4a", (53248 + 908) => x"00", (53248 + 909) => x"e0", (53248 + 910) => x"23", (53248 + 911) => x"d4", (53248 + 912) => x"60", (53248 + 913) => x"60", (53248 + 914) => x"f0", (53248 + 915) => x"18", (53248 + 916) => x"13", (53248 + 917) => x"94", (53248 + 918) => x"6e", (53248 + 919) => x"00", (53248 + 920) => x"13", (53248 + 921) => x"84", (53248 + 922) => x"41", (53248 + 923) => x"01", (53248 + 924) => x"74", (53248 + 925) => x"ff", (53248 + 926) => x"41", (53248 + 927) => x"04", (53248 + 928) => x"73", (53248 + 929) => x"ff", (53248 + 930) => x"41", (53248 + 931) => x"06", (53248 + 932) => x"73", (53248 + 933) => x"01", (53248 + 934) => x"41", (53248 + 935) => x"09", (53248 + 936) => x"74", (53248 + 937) => x"01", (53248 + 938) => x"00", (53248 + 939) => x"ee", (53248 + 940) => x"44", (53248 + 941) => x"00", (53248 + 942) => x"74", (53248 + 943) => x"01", (53248 + 944) => x"43", (53248 + 945) => x"00", (53248 + 946) => x"73", (53248 + 947) => x"01", (53248 + 948) => x"43", (53248 + 949) => x"38", (53248 + 950) => x"73", (53248 + 951) => x"ff", (53248 + 952) => x"44", (53248 + 953) => x"18", (53248 + 954) => x"74", (53248 + 955) => x"ff", (53248 + 956) => x"00", (53248 + 957) => x"ee", (53248 + 958) => x"6b", (53248 + 959) => x"00", (53248 + 960) => x"44", (53248 + 961) => x"00", (53248 + 962) => x"13", (53248 + 963) => x"ce", (53248 + 964) => x"43", (53248 + 965) => x"00", (53248 + 966) => x"13", (53248 + 967) => x"ce", (53248 + 968) => x"43", (53248 + 969) => x"3f", (53248 + 970) => x"13", (53248 + 971) => x"ce", (53248 + 972) => x"44", (53248 + 973) => x"1f", (53248 + 974) => x"6b", (53248 + 975) => x"bb", (53248 + 976) => x"6f", (53248 + 977) => x"00", (53248 + 978) => x"00", (53248 + 979) => x"ee", (53248 + 980) => x"63", (53248 + 981) => x"08", (53248 + 982) => x"64", (53248 + 983) => x"08", (53248 + 984) => x"a2", (53248 + 985) => x"29", (53248 + 986) => x"fe", (53248 + 987) => x"33", (53248 + 988) => x"f2", (53248 + 989) => x"65", (53248 + 990) => x"23", (53248 + 991) => x"ec", (53248 + 992) => x"63", (53248 + 993) => x"28", (53248 + 994) => x"a2", (53248 + 995) => x"29", (53248 + 996) => x"f6", (53248 + 997) => x"33", (53248 + 998) => x"f2", (53248 + 999) => x"65", (53248 + 1000) => x"23", (53248 + 1001) => x"f2", (53248 + 1002) => x"00", (53248 + 1003) => x"ee", (53248 + 1004) => x"f0", (53248 + 1005) => x"29", (53248 + 1006) => x"d3", (53248 + 1007) => x"45", (53248 + 1008) => x"73", (53248 + 1009) => x"06", (53248 + 1010) => x"f1", (53248 + 1011) => x"29", (53248 + 1012) => x"d3", (53248 + 1013) => x"45", (53248 + 1014) => x"73", (53248 + 1015) => x"06", (53248 + 1016) => x"f2", (53248 + 1017) => x"29", (53248 + 1018) => x"d3", (53248 + 1019) => x"45", (53248 + 1020) => x"00", (53248 + 1021) => x"ee", (53248 + 1022) => x"01", (53248 + 1023) => x"10", (53248 + 1024) => x"54", (53248 + 1025) => x"7c", (53248 + 1026) => x"6c", (53248 + 1027) => x"7c", (53248 + 1028) => x"7c", (53248 + 1029) => x"44", (53248 + 1030) => x"7c", (53248 + 1031) => x"7c", (53248 + 1032) => x"6c", (53248 + 1033) => x"7c", (53248 + 1034) => x"54", (53248 + 1035) => x"10", (53248 + 1036) => x"00", (53248 + 1037) => x"fc", (53248 + 1038) => x"78", (53248 + 1039) => x"6e", (53248 + 1040) => x"78", (53248 + 1041) => x"fc", (53248 + 1042) => x"00", (53248 + 1043) => x"3f", (53248 + 1044) => x"1e", (53248 + 1045) => x"76", (53248 + 1046) => x"1e", (53248 + 1047) => x"3f", (53248 + 1048) => x"00", (53248 + 1049) => x"80", (53248 + 1050) => x"a8", (53248 + 1051) => x"70", (53248 + 1052) => x"f8", (53248 + 1053) => x"70", (53248 + 1054) => x"a8", (53248 + 1055) => x"0b", (53248 + 1056) => x"1b", (53248 + 1057) => x"28", (53248 + 1058) => x"38", (53248 + 1059) => x"30", (53248 + 1060) => x"20", (53248 + 1061) => x"10", (53248 + 1062) => x"00", (53248 + 1063) => x"00", (53248 + 1064) => x"00", (53248 + 1065) => x"00", (53248 + 1066) => x"08", (53248 + 1067) => x"1b", (53248 + 1068) => x"1b", (53248 + 1069) => x"1b", (53248 + 1070) => x"18", (53248 + 1071) => x"04", 
                                
                                -- Vers by JMN
                                (57344 + 128) => x"03", (57344 + 129) => x"00", 
                                (57344 + 130) => x"00", (57344 + 131) => x"02",
                                (57344 + 132) => x"00", (57344 + 133) => x"1C",
                                (57344 + 134) => x"BF", (57344 + 135) => x"0E",
                                (57344 + 136) => x"00", (57344 + 137) => x"30", -- delay
                                (57344 + 138) => x"00",
                                (57344 + 512) => x"12", (57344 + 513) => x"1a", (57344 + 514) => x"4a", (57344 + 515) => x"4d", (57344 + 516) => x"4e", (57344 + 517) => x"20", (57344 + 518) => x"31", (57344 + 519) => x"39", (57344 + 520) => x"39", (57344 + 521) => x"31", (57344 + 522) => x"20", (57344 + 523) => x"53", (57344 + 524) => x"4f", (57344 + 525) => x"46", (57344 + 526) => x"54", (57344 + 527) => x"57", (57344 + 528) => x"41", (57344 + 529) => x"52", (57344 + 530) => x"45", (57344 + 531) => x"53", (57344 + 532) => x"20", (57344 + 533) => x"80", (57344 + 534) => x"80", (57344 + 535) => x"ff", (57344 + 536) => x"00", (57344 + 537) => x"00", (57344 + 538) => x"63", (57344 + 539) => x"00", (57344 + 540) => x"67", (57344 + 541) => x"00", (57344 + 542) => x"00", (57344 + 543) => x"e0", (57344 + 544) => x"a2", (57344 + 545) => x"17", (57344 + 546) => x"60", (57344 + 547) => x"00", (57344 + 548) => x"61", (57344 + 549) => x"00", (57344 + 550) => x"d0", (57344 + 551) => x"11", (57344 + 552) => x"71", (57344 + 553) => x"ff", (57344 + 554) => x"d0", (57344 + 555) => x"11", (57344 + 556) => x"71", (57344 + 557) => x"01", (57344 + 558) => x"70", (57344 + 559) => x"08", (57344 + 560) => x"30", (57344 + 561) => x"40", (57344 + 562) => x"12", (57344 + 563) => x"26", (57344 + 564) => x"71", (57344 + 565) => x"01", (57344 + 566) => x"a2", (57344 + 567) => x"15", (57344 + 568) => x"d0", (57344 + 569) => x"12", (57344 + 570) => x"70", (57344 + 571) => x"ff", (57344 + 572) => x"d0", (57344 + 573) => x"12", (57344 + 574) => x"70", (57344 + 575) => x"01", (57344 + 576) => x"71", (57344 + 577) => x"02", (57344 + 578) => x"31", (57344 + 579) => x"1f", (57344 + 580) => x"12", (57344 + 581) => x"38", (57344 + 582) => x"60", (57344 + 583) => x"08", (57344 + 584) => x"61", (57344 + 585) => x"10", (57344 + 586) => x"62", (57344 + 587) => x"04", (57344 + 588) => x"64", (57344 + 589) => x"37", (57344 + 590) => x"65", (57344 + 591) => x"0f", (57344 + 592) => x"66", (57344 + 593) => x"02", (57344 + 594) => x"d0", (57344 + 595) => x"11", (57344 + 596) => x"d4", (57344 + 597) => x"51", (57344 + 598) => x"68", (57344 + 599) => x"01", (57344 + 600) => x"e8", (57344 + 601) => x"a1", (57344 + 602) => x"62", (57344 + 603) => x"02", (57344 + 604) => x"68", (57344 + 605) => x"02", (57344 + 606) => x"e8", (57344 + 607) => x"a1", (57344 + 608) => x"62", (57344 + 609) => x"04", (57344 + 610) => x"68", (57344 + 611) => x"07", (57344 + 612) => x"e8", (57344 + 613) => x"a1", (57344 + 614) => x"62", (57344 + 615) => x"01", (57344 + 616) => x"68", (57344 + 617) => x"0a", (57344 + 618) => x"e8", (57344 + 619) => x"a1", (57344 + 620) => x"62", (57344 + 621) => x"03", (57344 + 622) => x"68", (57344 + 623) => x"0b", (57344 + 624) => x"e8", (57344 + 625) => x"a1", (57344 + 626) => x"66", (57344 + 627) => x"02", (57344 + 628) => x"68", (57344 + 629) => x"0f", (57344 + 630) => x"e8", (57344 + 631) => x"a1", (57344 + 632) => x"66", (57344 + 633) => x"04", (57344 + 634) => x"68", (57344 + 635) => x"0c", (57344 + 636) => x"e8", (57344 + 637) => x"a1", (57344 + 638) => x"66", (57344 + 639) => x"01", (57344 + 640) => x"68", (57344 + 641) => x"0d", (57344 + 642) => x"e8", (57344 + 643) => x"a1", (57344 + 644) => x"66", (57344 + 645) => x"03", (57344 + 646) => x"42", (57344 + 647) => x"01", (57344 + 648) => x"71", (57344 + 649) => x"ff", (57344 + 650) => x"42", (57344 + 651) => x"02", (57344 + 652) => x"70", (57344 + 653) => x"ff", (57344 + 654) => x"42", (57344 + 655) => x"03", (57344 + 656) => x"71", (57344 + 657) => x"01", (57344 + 658) => x"42", (57344 + 659) => x"04", (57344 + 660) => x"70", (57344 + 661) => x"01", (57344 + 662) => x"46", (57344 + 663) => x"01", (57344 + 664) => x"75", (57344 + 665) => x"ff", (57344 + 666) => x"46", (57344 + 667) => x"02", (57344 + 668) => x"74", (57344 + 669) => x"ff", (57344 + 670) => x"46", (57344 + 671) => x"03", (57344 + 672) => x"75", (57344 + 673) => x"01", (57344 + 674) => x"46", (57344 + 675) => x"04", (57344 + 676) => x"74", (57344 + 677) => x"01", (57344 + 678) => x"d0", (57344 + 679) => x"11", (57344 + 680) => x"3f", (57344 + 681) => x"00", (57344 + 682) => x"12", (57344 + 683) => x"b4", (57344 + 684) => x"d4", (57344 + 685) => x"51", (57344 + 686) => x"3f", (57344 + 687) => x"00", (57344 + 688) => x"12", (57344 + 689) => x"b8", (57344 + 690) => x"12", (57344 + 691) => x"56", (57344 + 692) => x"77", (57344 + 693) => x"01", (57344 + 694) => x"12", (57344 + 695) => x"ba", (57344 + 696) => x"73", (57344 + 697) => x"01", (57344 + 698) => x"68", (57344 + 699) => x"00", (57344 + 700) => x"78", (57344 + 701) => x"01", (57344 + 702) => x"38", (57344 + 703) => x"00", (57344 + 704) => x"12", (57344 + 705) => x"bc", (57344 + 706) => x"00", (57344 + 707) => x"e0", (57344 + 708) => x"60", (57344 + 709) => x"08", (57344 + 710) => x"61", (57344 + 711) => x"04", (57344 + 712) => x"f3", (57344 + 713) => x"29", (57344 + 714) => x"d0", (57344 + 715) => x"15", (57344 + 716) => x"60", (57344 + 717) => x"34", (57344 + 718) => x"f7", (57344 + 719) => x"29", (57344 + 720) => x"d0", (57344 + 721) => x"15", (57344 + 722) => x"68", (57344 + 723) => x"00", (57344 + 724) => x"78", (57344 + 725) => x"01", (57344 + 726) => x"38", (57344 + 727) => x"00", (57344 + 728) => x"12", (57344 + 729) => x"d4", (57344 + 730) => x"43", (57344 + 731) => x"08", (57344 + 732) => x"12", (57344 + 733) => x"e4", (57344 + 734) => x"47", (57344 + 735) => x"08", (57344 + 736) => x"12", (57344 + 737) => x"e4", (57344 + 738) => x"12", (57344 + 739) => x"1e", (57344 + 740) => x"12", (57344 + 741) => x"e4", 
                                others => ( others => '0')
                            );
    signal read_address : std_logic_vector( 15 downto 0 );
begin

    process ( clock )
    begin
        if ( rising_edge( clock ) ) then
            if( we = '1' ) then
                sys_RAM( to_integer( unsigned( address ))) <= dataIn;
            end if;
            
            read_address <= address;
        end if;
    end process;

    dataOut <= sys_RAM( to_integer( unsigned( read_address )));
end Behavioral;
